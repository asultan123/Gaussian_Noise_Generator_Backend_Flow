* Nettran: AMD.64 Release B-2008.09.SP5.26004 2012/07/19
* Created:  4/21/2018  15:58
* Options: -rootCell gng -verilog-b0 VSS -verilog-b1 VDD -sp /home/standard_cell_libraries/NangateOpenCellLibrary_PDKv1_3_v2010_12/lib/Back_End/spice/NangateOpenCellLibrary.spi -verilog /home/mohamed/Desktop/ref_flow/pnr/output_verilog_withphysical -outType spice -outName gng.sp 

.GLOBAL VDD VSS 

.SUBCKT XOR2_X2 A B Z VDD VSS 
M_i_41_29 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47_27 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_18 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_35 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19_23 net_001b A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24_4 VSS B net_001b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XNOR2_X2 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_25 VDD B net_003b VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48_8 net_003b A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42_14 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_23_12 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17_20 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11_23 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT TLAT_X1 D G OE Q VDD VSS 
M_i_111 Q net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_106 net_010 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_91 net_005 OE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_99 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 VDD net_006 net_009 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_81 net_009 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_003 net_000 net_008 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_70 net_008 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_64 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 Q OE net_007 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_47 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_34 net_005 OE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TINV_X1 EN I ZN VDD VSS 
M_i_29 ZN EN net_002 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24 net_002 I VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VDD EN net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 ZN net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_7 net_001 I VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0 VSS EN net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TBUF_X8 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X4 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X2 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X16 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_10 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_83 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_42 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_51 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9_17 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18_103 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39_66 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50_12 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_116 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_106 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_120 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_43 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42_108 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37_112 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45_122 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40_125 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X1 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT SDFF_X2 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_115_2 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108_51 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7_4 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_50 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFF_X1 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFS_X2 D SE SI SN CK Q QN VDD VSS 
M_i_230_17 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237_1 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103_26 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110_2 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 VSS net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_93 net_014 SN net_015 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFS_X1 D SE SI SN CK Q QN VDD VSS 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 net_015 net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_93 net_014 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFR_X2 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_116_1 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123_146 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_10 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7_145 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFR_X1 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X2 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_277_67 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290_11 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 net_013 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_106 net_017 SN net_016 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_119 net_019 RN net_018 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_114 net_018 net_017 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_125_68 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132_2 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X1 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_106 net_017 net_013 net_016 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_114 net_018 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_119 net_019 net_017 net_018 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 ZN_neg A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT OR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_1__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m0 VDD A2 net_0__m0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m0 net_0__m0_0__m0_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m1 ZN_neg A1 net_0__m0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m1 net_0__m0_0__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 ZN VDD VSS 
M_i_8 VDD A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 B3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 ZN A3 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_0 B3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 VDD A2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_1__m3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN A1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_1__m2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 VDD B2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 net_2__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN B1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 net_2__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_1 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_0 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_5 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 A1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_0 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_1 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_5 A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 ZN A1 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A2 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 ZN C1 net_4__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 net_4__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 VDD C2 net_4__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 net_4__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0__m1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_3_x4_0 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_1 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_2 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_3 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN_4 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_4 C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_7_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 VDD B2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 net_1__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN B1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_1__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X4 A B C1 C2 ZN VDD VSS 
M_i_5__m3 VDD C2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_2__m3 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN C1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_2__m2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_0 A net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_1__m3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7_1_96 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_102 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34_44 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_56 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_88 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24_95 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_68 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6_75 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8_108 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_109 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_8 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29_45 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_52 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_79 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13_89 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_77 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22_71 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5_83 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_65 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_56 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_52 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_43 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_34 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_24 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_85 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_67 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_58 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_49 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_40 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_31 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5_1_m2__m1 VDD A3 net_1_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m1 net_1_0__m1 A2 net_0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m1 net_0_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m0 ZN A1 net_0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m0 net_0_0__m0_0 A2 net_1_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1_m2__m0 net_1_0__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0_x2__m1 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m1 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m0 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2__m0 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_52 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_154 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_49 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_100 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_202 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_87 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_36 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_189 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_15 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_66 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_168 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_17 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_68 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_170 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_43 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_94 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_196 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_75 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_24 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_177 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_34 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_85 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_187 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5__m3 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m3 VSS A3 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m3 net_1__m3 A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5__m0_x2__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_2__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_x2__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m1 VSS A2 net_0__m0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X2 A B S Z VDD VSS 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_1_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 Z_neg B net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_2 x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS x1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT LOGIC1_X1 Z VDD VSS 
M_p_tran_2 VDD A Z VDD PMOS_VTL L=0.050000U W=0.135000U 
M_n_tran_1 VSS A A VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT FILLCELL_X8 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X4 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X32 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X2 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X16 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X1 VDD VSS 
.ENDS

.SUBCKT DLL_X2 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_92_11 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_42_3 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLL_X1 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X2 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_89 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_41 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X1 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X2 D SN CK Q QN VDD VSS 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189_10 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182_20 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86_15 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79_29 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X1 D SN CK Q QN VDD VSS 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X2 D RN CK Q QN VDD VSS 
M_i_187_39 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180_3 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83_49 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76_4 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X1 D RN CK Q QN VDD VSS 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFRS_X2 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP81_1_55 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0_51 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 z41 z56 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN51 VSS RN nn5 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN91_0_0_58 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81_53 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFFRS_X1 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 RN z56 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN51 VSS z41 nn5 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X8 CK E GCK VDD VSS 
M_i_109_4_19_36 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24_52 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_22 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_53 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74_97 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71_87 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_99 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_72 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57_165 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7_25_30 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10_28 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_58 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_40 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66_78 VSS net_000 net_007d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75_82 net_007d CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_71 net_007c CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_63 VSS net_000 net_007c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_174 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X4 CK E GCK VDD VSS 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X2 CK E GCK VDD VSS 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X1 CK E GCK VDD VSS 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X8 CK E SE GCK VDD VSS 
M_i_133_10_28_7 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11_14 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_20 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_38 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72_145 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69_164 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_158 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_163 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101_94 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29_4 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15_27 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_55 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_12 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76_137 net_008d CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77_169 net_007 net_002 net_008d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_123 net_007 net_002 net_008c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_150 net_008c CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33_93 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X4 CK E SE GCK VDD VSS 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X2 CK E SE GCK VDD VSS 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X1 CK E SE GCK VDD VSS 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT BUF_X8 A Z VDD VSS 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X4 A Z VDD VSS 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 VSS B2 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_1__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 ZN B1 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 net_1__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_0 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_1 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A2 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_5 A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_1 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_0 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 C1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_5 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_7__m0 net_3 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0 net_0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_2__m0_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN C1 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_2__m1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_0_x4_3 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_2 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_1 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_0 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN_4 C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_4 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 net_2 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS B2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN B1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS B2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN B1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m0_x2__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m0 VSS B2 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 net_0__m0_0__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 ZN B1 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_0__m0_0__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X4 A B C1 C2 ZN VDD VSS 
M_i_11_3 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_2 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_0 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_1 VDD ZN_3 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_0 ZN_4 ZN_3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 C2 ZN_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_3 C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10_3 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_2 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_1 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_1 VSS ZN_3 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_0 ZN_4 ZN_3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 net_1 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1 B net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT ANTENNA_X1 A VDD VSS 
.ENDS

.SUBCKT AND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 x1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A2 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 x1 A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A1 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 x1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 VDD A3 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 x1 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0__m1 A1 x1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 x1 A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_0_x4_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m1 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m0 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_4__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 VSS A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X4 A1 A2 ZN VDD VSS 
M_i_2_3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_3 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_2 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_0 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X4 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m1_58 VDD A2 net_0__m0__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1_45 net_0__m0__m2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0_52 ZN A1 net_0__m0__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0_38 net_0__m0__m3 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m1_23 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1_57 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0_35 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0_16 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFF_X2 D CK Q QN VDD VSS 
M_MP13_26 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14_5 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13_38 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14_8 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKBUF_X3 A Z VDD VSS 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN C1 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_2 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 ZN C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NOR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X2 A Z VDD VSS 
M_i_1_0_x2_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X1 A B S Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B net_3 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_3 x1 Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_5 Z_neg x1 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_1 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 VDD A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X16 A Z VDD VSS 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X2 A ZN VDD VSS 
M_i_1_0_x2_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT LOGIC0_X1 Z VDD VSS 
M_transistor_0 VDD A A VDD PMOS_VTL L=0.050000U W=0.090000U 
M_n_tran_1 VSS A Z VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT DFF_X1 D CK Q QN VDD VSS 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKBUF_X2 A Z VDD VSS 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT XNOR2_X1 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NOR2_X1 A1 A2 ZN VDD VSS 
M_i_2 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X1 A1 A2 ZN VDD VSS 
M_i_2 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XOR2_X1 A B Z VDD VSS 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AND2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT INV_X4 A ZN VDD VSS 
M_i_1_0_x4_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X8 A ZN VDD VSS 
M_i_1_0_x8_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x8_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X32 A Z VDD VSS 
M_i_1_31 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_14 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_13 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_12 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_11 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_10 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_9 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_15 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_14 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_13 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_12 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_11 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_10 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_9 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_8 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT HA_X1 A B CO S VDD VSS 
M_i_11 CO CO_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15 VDD B CO_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_14 CO_neg A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 x1 A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_2 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD x1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 A S VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 S B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 CO CO_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS B net_3 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_12 net_3 A CO_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_6 VSS A x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 x1 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS x1 S VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 S A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VSS B net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X1 A ZN VDD VSS 
M_i_1 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT FA_X1 A B CI CO S VDD VSS 
M_instance_315 S net_005 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_275 VDD A net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_280 net_009 B net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_284 net_010 CI net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_290 net_005 net_001 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_303 net_011 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_297 VDD CI net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_309 net_011 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_263 VDD B net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_269 net_008 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_257 net_001 CI net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_251 net_007 A net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_246 VDD B net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_239 CO net_001 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_233 S net_005 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_instance_194 VSS A net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_199 net_003 B net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_203 net_004 CI net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_209 net_005 net_001 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_221 net_006 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_215 VSS CI net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_227 net_006 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_182 VSS B net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_188 net_002 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_176 net_001 CI net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_170 net_000 A net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_166 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_159 CO net_001 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X16 A ZN VDD VSS 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKBUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.095000U 
.ENDS

.SUBCKT BUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT INV_X32 A ZN VDD VSS 
M_i_1_31 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT gng_lzd data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] 
+ data_in[60] data_in[59] data_in[58] data_in[57] data_in[56] data_in[55] data_in[54] 
+ data_in[53] data_in[52] data_in[51] data_in[50] data_in[49] data_in[48] data_in[47] 
+ data_in[46] data_in[45] data_in[44] data_in[43] data_in[42] data_in[41] data_in[40] 
+ data_in[39] data_in[38] data_in[37] data_in[36] data_in[35] data_in[34] data_in[33] 
+ data_in[32] data_in[31] data_in[30] data_in[29] data_in[28] data_in[27] data_in[26] 
+ data_in[25] data_in[24] data_in[23] data_in[22] data_in[21] data_in[20] data_in[19] 
+ data_in[18] data_in[17] data_in[16] data_in[15] data_in[14] data_in[13] data_in[12] 
+ data_in[11] data_in[10] data_in[9] data_in[8] data_in[7] data_in[6] data_in[5] 
+ data_in[4] data_in[3] data_in[2] data_in[1] data_in[0] 
XU22 n58 n15 n18 n14 n56 NETTRAN_DUMMY_1 NETTRAN_DUMMY_2 OAI22_X1 
XU21 n54 n34 n33 n39 n51 NETTRAN_DUMMY_3 NETTRAN_DUMMY_4 OAI22_X1 
XU20 n45 n5 NETTRAN_DUMMY_5 NETTRAN_DUMMY_6 INV_X1 
XU19 n48 n22 NETTRAN_DUMMY_7 NETTRAN_DUMMY_8 INV_X1 
XU18 data_out[5] n48 n43 NETTRAN_DUMMY_9 NETTRAN_DUMMY_10 NAND2_X1 
XU17 n55 n2 NETTRAN_DUMMY_11 NETTRAN_DUMMY_12 INV_X1 
XU16 n55 n130 n42 NETTRAN_DUMMY_13 NETTRAN_DUMMY_14 NAND2_X1 
XU15 n42 n43 data_out[4] NETTRAN_DUMMY_15 NETTRAN_DUMMY_16 NAND2_X1 
XU14 n55 n56 n57 n2 n49 NETTRAN_DUMMY_17 NETTRAN_DUMMY_18 AOI22_X1 
XU13 n48 n51 n52 n22 n50 NETTRAN_DUMMY_19 NETTRAN_DUMMY_20 AOI22_X1 
XU12 data_out[5] n49 n50 n130 n134 NETTRAN_DUMMY_21 NETTRAN_DUMMY_22 OAI22_X1 
XU11 n130 n48 n24 n46 NETTRAN_DUMMY_23 NETTRAN_DUMMY_24 NOR3_X1 
XU10 n46 n45 n2 n44 NETTRAN_DUMMY_25 NETTRAN_DUMMY_26 AOI21_X1 
XU9 n44 n33 n43 n14 n42 n131 NETTRAN_DUMMY_27 NETTRAN_DUMMY_28 OAI221_X1 
XU8 n55 n70 n71 n2 n59 NETTRAN_DUMMY_29 NETTRAN_DUMMY_30 AOI22_X1 
XU7 n67 n37 n68 n35 n69 n40 n60 NETTRAN_DUMMY_31 NETTRAN_DUMMY_32 AOI222_X1 
XU6 n61 data_out[5] n59 n60 n43 n133 NETTRAN_DUMMY_33 NETTRAN_DUMMY_34 OAI221_X1 
XU5 n91 n92 n93 n94 n83 NETTRAN_DUMMY_35 NETTRAN_DUMMY_36 NOR4_X1 
XU4 n85 n86 n87 n88 n84 NETTRAN_DUMMY_37 NETTRAN_DUMMY_38 NOR4_X1 
XU3 n82 n130 n55 n83 n84 n42 n132 NETTRAN_DUMMY_39 NETTRAN_DUMMY_40 OAI222_X1 
XU2 data_in[55] data_in[56] data_in[54] n98 n45 NETTRAN_DUMMY_41 NETTRAN_DUMMY_42 NOR4_X1 
XU76 data_in[13] n23 data_in[15] data_in[14] n48 NETTRAN_DUMMY_43 NETTRAN_DUMMY_44 NOR4_X1 
XU44 data_in[45] n4 data_in[47] data_in[46] n55 NETTRAN_DUMMY_45 NETTRAN_DUMMY_46 NOR4_X2 
XU117 data_in[47] n11 NETTRAN_DUMMY_47 NETTRAN_DUMMY_48 INV_X1 
XU116 data_in[35] n19 NETTRAN_DUMMY_49 NETTRAN_DUMMY_50 INV_X1 
XU115 data_in[51] n10 NETTRAN_DUMMY_51 NETTRAN_DUMMY_52 INV_X1 
XU114 n89 data_in[44] n78 NETTRAN_DUMMY_53 NETTRAN_DUMMY_54 OR2_X1 
XU113 n95 data_in[60] n73 NETTRAN_DUMMY_55 NETTRAN_DUMMY_56 OR2_X1 
XU112 data_in[26] n27 NETTRAN_DUMMY_57 NETTRAN_DUMMY_58 INV_X1 
XU111 n64 data_in[27] n27 n102 NETTRAN_DUMMY_59 NETTRAN_DUMMY_60 OAI21_X1 
XU110 data_in[43] n16 NETTRAN_DUMMY_61 NETTRAN_DUMMY_62 INV_X1 
XU109 n78 data_in[42] n16 n88 NETTRAN_DUMMY_63 NETTRAN_DUMMY_64 AOI21_X1 
XU108 data_in[59] n7 NETTRAN_DUMMY_65 NETTRAN_DUMMY_66 INV_X1 
XU107 n73 data_in[58] n7 n94 NETTRAN_DUMMY_67 NETTRAN_DUMMY_68 AOI21_X1 
XU106 n114 data_in[12] n68 NETTRAN_DUMMY_69 NETTRAN_DUMMY_70 NOR2_X1 
XU105 n108 data_in[28] n64 NETTRAN_DUMMY_71 NETTRAN_DUMMY_72 NOR2_X1 
XU104 data_in[2] data_in[1] data_in[4] data_in[3] n113 NETTRAN_DUMMY_73 NETTRAN_DUMMY_74 NOR4_X1 
XU103 data_in[37] n15 n99 NETTRAN_DUMMY_75 NETTRAN_DUMMY_76 OR2_X1 
XU102 data_in[39] data_in[40] data_in[38] n99 n58 NETTRAN_DUMMY_77 NETTRAN_DUMMY_78 NOR4_X1 
XU101 data_in[23] n28 NETTRAN_DUMMY_79 NETTRAN_DUMMY_80 INV_X1 
XU100 data_in[27] n26 NETTRAN_DUMMY_81 NETTRAN_DUMMY_82 INV_X1 
XU99 n65 n28 n63 n26 n64 n62 NETTRAN_DUMMY_83 NETTRAN_DUMMY_84 AOI221_X1 
XU98 n62 n48 n130 n61 NETTRAN_DUMMY_85 NETTRAN_DUMMY_86 OR3_X1 
XU97 data_in[0] n33 n39 n112 NETTRAN_DUMMY_87 NETTRAN_DUMMY_88 OR3_X1 
XU96 n58 data_in[40] n15 n77 NETTRAN_DUMMY_89 NETTRAN_DUMMY_90 OR3_X1 
XU95 n45 data_in[56] n6 n72 NETTRAN_DUMMY_91 NETTRAN_DUMMY_92 OR3_X1 
XU94 data_in[6] n38 NETTRAN_DUMMY_93 NETTRAN_DUMMY_94 INV_X1 
XU93 n67 data_in[7] n38 n109 NETTRAN_DUMMY_95 NETTRAN_DUMMY_96 OAI21_X1 
XU92 data_in[22] n29 NETTRAN_DUMMY_97 NETTRAN_DUMMY_98 INV_X1 
XU91 n63 data_in[23] n29 n103 NETTRAN_DUMMY_99 NETTRAN_DUMMY_100 OAI21_X1 
XU90 data_in[2] n41 NETTRAN_DUMMY_101 NETTRAN_DUMMY_102 INV_X1 
XU89 n69 data_in[3] n41 n110 NETTRAN_DUMMY_103 NETTRAN_DUMMY_104 OAI21_X1 
XU88 data_in[18] n31 NETTRAN_DUMMY_105 NETTRAN_DUMMY_106 INV_X1 
XU87 n66 data_in[19] n31 n104 NETTRAN_DUMMY_107 NETTRAN_DUMMY_108 OAI21_X1 
XU86 data_in[14] n32 NETTRAN_DUMMY_109 NETTRAN_DUMMY_110 INV_X1 
XU85 n106 data_in[15] n32 n105 NETTRAN_DUMMY_111 NETTRAN_DUMMY_112 OAI21_X1 
XU84 n80 n13 NETTRAN_DUMMY_113 NETTRAN_DUMMY_114 INV_X1 
XU83 n13 data_in[30] n20 n85 NETTRAN_DUMMY_115 NETTRAN_DUMMY_116 AOI21_X1 
XU82 n4 data_in[46] n11 n91 NETTRAN_DUMMY_117 NETTRAN_DUMMY_118 AOI21_X1 
XU81 n81 n12 NETTRAN_DUMMY_119 NETTRAN_DUMMY_120 INV_X1 
XU80 n12 data_in[34] n19 n86 NETTRAN_DUMMY_121 NETTRAN_DUMMY_122 AOI21_X1 
XU79 n76 n1 NETTRAN_DUMMY_123 NETTRAN_DUMMY_124 INV_X1 
XU78 n1 data_in[50] n10 n92 NETTRAN_DUMMY_125 NETTRAN_DUMMY_126 AOI21_X1 
XU77 data_in[39] n17 NETTRAN_DUMMY_127 NETTRAN_DUMMY_128 INV_X1 
XU75 n77 data_in[38] n17 n87 NETTRAN_DUMMY_129 NETTRAN_DUMMY_130 AOI21_X1 
XU74 data_in[55] n8 NETTRAN_DUMMY_131 NETTRAN_DUMMY_132 INV_X1 
XU73 n72 data_in[54] n8 n93 NETTRAN_DUMMY_133 NETTRAN_DUMMY_134 AOI21_X1 
XU72 n66 n21 NETTRAN_DUMMY_135 NETTRAN_DUMMY_136 INV_X1 
XU71 n23 data_in[15] n21 data_in[19] n65 NETTRAN_DUMMY_137 NETTRAN_DUMMY_138 OAI22_X1 
XU70 n75 n11 n76 n10 n74 NETTRAN_DUMMY_139 NETTRAN_DUMMY_140 AOI22_X1 
XU69 n74 data_in[55] n72 data_in[59] n73 n71 NETTRAN_DUMMY_141 NETTRAN_DUMMY_142 OAI221_X1 
XU68 n80 n20 n81 n19 n79 NETTRAN_DUMMY_143 NETTRAN_DUMMY_144 AOI22_X1 
XU67 n79 data_in[39] n77 data_in[43] n78 n70 NETTRAN_DUMMY_145 NETTRAN_DUMMY_146 OAI221_X1 
XU66 n68 data_in[11] n36 n111 NETTRAN_DUMMY_147 NETTRAN_DUMMY_148 OAI21_X1 
XU65 n102 n103 n104 n105 n101 NETTRAN_DUMMY_149 NETTRAN_DUMMY_150 NAND4_X1 
XU64 n109 n110 n111 n112 n100 NETTRAN_DUMMY_151 NETTRAN_DUMMY_152 NAND4_X1 
XU63 n48 n100 n101 n22 n82 NETTRAN_DUMMY_153 NETTRAN_DUMMY_154 AOI22_X1 
XU62 n113 data_in[4] n33 n69 NETTRAN_DUMMY_155 NETTRAN_DUMMY_156 NOR3_X1 
XU61 n90 data_in[36] n14 n81 NETTRAN_DUMMY_157 NETTRAN_DUMMY_158 NOR3_X1 
XU60 n96 data_in[52] n5 n76 NETTRAN_DUMMY_159 NETTRAN_DUMMY_160 NOR3_X1 
XU59 n54 data_in[8] n34 n67 NETTRAN_DUMMY_161 NETTRAN_DUMMY_162 NOR3_X1 
XU58 n53 data_in[24] n25 n63 NETTRAN_DUMMY_163 NETTRAN_DUMMY_164 NOR3_X1 
XU57 n107 data_in[20] n24 n66 NETTRAN_DUMMY_165 NETTRAN_DUMMY_166 NOR3_X1 
XU56 data_in[16] n30 n24 n106 NETTRAN_DUMMY_167 NETTRAN_DUMMY_168 NOR3_X1 
XU55 data_in[48] n9 n5 n75 NETTRAN_DUMMY_169 NETTRAN_DUMMY_170 NOR3_X1 
XU54 data_in[58] data_in[57] data_in[60] data_in[59] n95 NETTRAN_DUMMY_171 NETTRAN_DUMMY_172 NOR4_X1 
XU53 data_in[42] data_in[41] data_in[44] data_in[43] n89 NETTRAN_DUMMY_173 NETTRAN_DUMMY_174 NOR4_X1 
XU52 data_in[32] n18 n14 n80 NETTRAN_DUMMY_175 NETTRAN_DUMMY_176 NOR3_X1 
XU51 data_in[29] data_in[31] data_in[30] n97 NETTRAN_DUMMY_177 NETTRAN_DUMMY_178 NOR3_X1 
XU50 n80 n55 n97 n47 NETTRAN_DUMMY_179 NETTRAN_DUMMY_180 NAND3_X1 
XU49 data_in[26] data_in[25] data_in[28] data_in[27] n108 NETTRAN_DUMMY_181 NETTRAN_DUMMY_182 NOR4_X1 
XU48 data_in[11] data_in[10] data_in[9] data_in[12] n114 NETTRAN_DUMMY_183 NETTRAN_DUMMY_184 NOR4_X1 
XU47 data_in[34] data_in[33] data_in[36] data_in[35] n90 NETTRAN_DUMMY_185 NETTRAN_DUMMY_186 NOR4_X1 
XU46 data_in[50] data_in[49] data_in[52] data_in[51] n96 NETTRAN_DUMMY_187 NETTRAN_DUMMY_188 NOR4_X1 
XU45 data_in[18] data_in[17] data_in[20] data_in[19] n107 NETTRAN_DUMMY_189 NETTRAN_DUMMY_190 NOR4_X1 
XU43 data_in[21] n25 n116 NETTRAN_DUMMY_191 NETTRAN_DUMMY_192 OR2_X1 
XU42 data_in[23] data_in[24] data_in[22] n116 n53 NETTRAN_DUMMY_193 NETTRAN_DUMMY_194 NOR4_X1 
XU41 data_in[5] n34 n115 NETTRAN_DUMMY_195 NETTRAN_DUMMY_196 OR2_X1 
XU40 data_in[7] data_in[8] data_in[6] n115 n54 NETTRAN_DUMMY_197 NETTRAN_DUMMY_198 NOR4_X1 
XU39 data_in[53] n6 n98 NETTRAN_DUMMY_199 NETTRAN_DUMMY_200 OR2_X1 
XU38 n113 n39 NETTRAN_DUMMY_201 NETTRAN_DUMMY_202 INV_X1 
XU37 n75 n4 NETTRAN_DUMMY_203 NETTRAN_DUMMY_204 INV_X1 
XU36 n106 n23 NETTRAN_DUMMY_205 NETTRAN_DUMMY_206 INV_X1 
XU35 n90 n18 NETTRAN_DUMMY_207 NETTRAN_DUMMY_208 INV_X1 
XU34 n96 n9 NETTRAN_DUMMY_209 NETTRAN_DUMMY_210 INV_X1 
XU33 n107 n30 NETTRAN_DUMMY_211 NETTRAN_DUMMY_212 INV_X1 
XU32 n95 n6 NETTRAN_DUMMY_213 NETTRAN_DUMMY_214 INV_X1 
XU31 n89 n15 NETTRAN_DUMMY_215 NETTRAN_DUMMY_216 INV_X1 
XU30 n108 n25 NETTRAN_DUMMY_217 NETTRAN_DUMMY_218 INV_X1 
XU29 n114 n34 NETTRAN_DUMMY_219 NETTRAN_DUMMY_220 INV_X1 
XU28 n130 data_out[5] NETTRAN_DUMMY_221 NETTRAN_DUMMY_222 INV_X1 
XU27 n53 n25 n30 n24 n52 NETTRAN_DUMMY_223 NETTRAN_DUMMY_224 OAI22_X1 
XU26 n45 n6 n9 n5 n57 NETTRAN_DUMMY_225 NETTRAN_DUMMY_226 OAI22_X1 
XU25 n58 n14 NETTRAN_DUMMY_227 NETTRAN_DUMMY_228 INV_X1 
XU24 n54 n33 NETTRAN_DUMMY_229 NETTRAN_DUMMY_230 INV_X1 
XU23 n53 n24 NETTRAN_DUMMY_231 NETTRAN_DUMMY_232 INV_X1 
XU122 data_in[10] n36 NETTRAN_DUMMY_233 NETTRAN_DUMMY_234 INV_X1 
XU121 data_in[7] n37 NETTRAN_DUMMY_235 NETTRAN_DUMMY_236 INV_X1 
XU120 data_in[11] n35 NETTRAN_DUMMY_237 NETTRAN_DUMMY_238 INV_X1 
XU119 data_in[3] n40 NETTRAN_DUMMY_239 NETTRAN_DUMMY_240 INV_X1 
XU118 data_in[31] n20 NETTRAN_DUMMY_241 NETTRAN_DUMMY_242 INV_X1 
XU1 n131 n3 NETTRAN_DUMMY_243 NETTRAN_DUMMY_244 INV_X1 
XU123 n3 data_out[3] NETTRAN_DUMMY_245 NETTRAN_DUMMY_246 INV_X32 
XU124 n134 n118 NETTRAN_DUMMY_247 NETTRAN_DUMMY_248 INV_X1 
XU125 n118 n119 NETTRAN_DUMMY_249 NETTRAN_DUMMY_250 INV_X32 
XU126 n119 n120 NETTRAN_DUMMY_251 NETTRAN_DUMMY_252 INV_X1 
XU127 n120 data_out[2] NETTRAN_DUMMY_253 NETTRAN_DUMMY_254 INV_X32 
XU128 n133 n122 NETTRAN_DUMMY_255 NETTRAN_DUMMY_256 INV_X1 
XU129 n122 n123 NETTRAN_DUMMY_257 NETTRAN_DUMMY_258 INV_X32 
XU130 n123 n124 NETTRAN_DUMMY_259 NETTRAN_DUMMY_260 INV_X1 
XU131 n124 data_out[1] NETTRAN_DUMMY_261 NETTRAN_DUMMY_262 INV_X32 
XU132 n127 n126 NETTRAN_DUMMY_263 NETTRAN_DUMMY_264 CLKBUF_X1 
XU133 n132 n127 NETTRAN_DUMMY_265 NETTRAN_DUMMY_266 INV_X1 
XU134 n126 data_out[0] NETTRAN_DUMMY_267 NETTRAN_DUMMY_268 INV_X32 
XU135 n47 n129 NETTRAN_DUMMY_269 NETTRAN_DUMMY_270 INV_X32 
XU136 n129 n130 NETTRAN_DUMMY_271 NETTRAN_DUMMY_272 INV_X1 
.ENDS

.SUBCKT gng_coef c2[16] c2[15] c2[14] c2[13] c2[12] c2[11] c2[10] c2[9] c2[8] c2[7] 
+ c2[6] c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] clk c1[17] c1[16] c1[15] c1[14] c1[13] 
+ c1[12] c1[11] c1[10] c1[9] c1[8] c1[7] c1[6] c1[5] c1[4] c1[3] c1[2] c1[1] c1[0] 
+ c0[17] c0[16] c0[15] c0[14] c0[13] c0[12] c0[11] c0[10] c0[9] c0[8] c0[7] c0[6] 
+ c0[5] c0[4] c0[3] c0[2] c0[1] c0[0] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] 
+ addr[1] addr[0] IN0 IN1 IN2 IN3 IN4 IN5 clk_cts_0 clk_cts_1 
XU1834 n488 n492 n1547 NETTRAN_DUMMY_273 NETTRAN_DUMMY_274 XOR2_X1 
XU1832 n537 n1545 NETTRAN_DUMMY_275 NETTRAN_DUMMY_276 INV_X1 
XU1831 n548 n1544 NETTRAN_DUMMY_277 NETTRAN_DUMMY_278 INV_X1 
XU1830 n539 n1543 NETTRAN_DUMMY_279 NETTRAN_DUMMY_280 INV_X1 
XU1829 n601 n1542 NETTRAN_DUMMY_281 NETTRAN_DUMMY_282 INV_X1 
XU1828 n627 n1541 NETTRAN_DUMMY_283 NETTRAN_DUMMY_284 INV_X1 
XU1827 n6 n1540 NETTRAN_DUMMY_285 NETTRAN_DUMMY_286 INV_X1 
XU1826 n525 n1539 NETTRAN_DUMMY_287 NETTRAN_DUMMY_288 INV_X1 
XU1825 n536 n1538 NETTRAN_DUMMY_289 NETTRAN_DUMMY_290 INV_X1 
XU1824 n1 n1537 NETTRAN_DUMMY_291 NETTRAN_DUMMY_292 INV_X1 
XU1637 addr[0] n515 NETTRAN_DUMMY_293 NETTRAN_DUMMY_294 BUF_X2 
XU1635 addr[0] n513 NETTRAN_DUMMY_295 NETTRAN_DUMMY_296 BUF_X1 
XU1631 addr[0] n509 NETTRAN_DUMMY_297 NETTRAN_DUMMY_298 BUF_X2 
XU1629 addr[1] n507 NETTRAN_DUMMY_299 NETTRAN_DUMMY_300 BUF_X2 
XU1625 addr[1] n503 NETTRAN_DUMMY_301 NETTRAN_DUMMY_302 BUF_X2 
XU1624 addr[1] n502 NETTRAN_DUMMY_303 NETTRAN_DUMMY_304 BUF_X2 
XU1622 addr[1] n500 NETTRAN_DUMMY_305 NETTRAN_DUMMY_306 BUF_X2 
XU1621 addr[1] n499 NETTRAN_DUMMY_307 NETTRAN_DUMMY_308 BUF_X2 
XU1619 addr[1] n497 NETTRAN_DUMMY_309 NETTRAN_DUMMY_310 BUF_X1 
XU1617 addr[1] n495 NETTRAN_DUMMY_311 NETTRAN_DUMMY_312 BUF_X1 
XU1615 IN0 n492 NETTRAN_DUMMY_313 NETTRAN_DUMMY_314 CLKBUF_X2 
XU1597 IN1 n487 NETTRAN_DUMMY_315 NETTRAN_DUMMY_316 BUF_X2 
XU1595 IN1 n484 NETTRAN_DUMMY_317 NETTRAN_DUMMY_318 BUF_X2 
XU1591 IN1 n480 NETTRAN_DUMMY_319 NETTRAN_DUMMY_320 BUF_X2 
XU822 IN2 n477 NETTRAN_DUMMY_321 NETTRAN_DUMMY_322 BUF_X2 
XU707 IN2 n475 NETTRAN_DUMMY_323 NETTRAN_DUMMY_324 BUF_X2 
XU568 IN2 n473 NETTRAN_DUMMY_325 NETTRAN_DUMMY_326 BUF_X2 
XU534 IN2 n471 NETTRAN_DUMMY_327 NETTRAN_DUMMY_328 BUF_X1 
XU521 IN2 n468 NETTRAN_DUMMY_329 NETTRAN_DUMMY_330 BUF_X1 
XU504 IN2 n466 NETTRAN_DUMMY_331 NETTRAN_DUMMY_332 BUF_X2 
XU497 IN2 n464 NETTRAN_DUMMY_333 NETTRAN_DUMMY_334 BUF_X2 
XU491 IN2 n462 NETTRAN_DUMMY_335 NETTRAN_DUMMY_336 BUF_X2 
XU486 IN2 n460 NETTRAN_DUMMY_337 NETTRAN_DUMMY_338 BUF_X2 
XU484 IN2 n458 NETTRAN_DUMMY_339 NETTRAN_DUMMY_340 BUF_X2 
XU481 IN3 n455 NETTRAN_DUMMY_341 NETTRAN_DUMMY_342 BUF_X1 
XU259 IN3 n454 NETTRAN_DUMMY_343 NETTRAN_DUMMY_344 BUF_X2 
XU201 IN3 n453 NETTRAN_DUMMY_345 NETTRAN_DUMMY_346 BUF_X2 
XU147 IN3 n452 NETTRAN_DUMMY_347 NETTRAN_DUMMY_348 BUF_X2 
XU49 IN3 n448 NETTRAN_DUMMY_349 NETTRAN_DUMMY_350 BUF_X2 
XU46 IN4 n445 NETTRAN_DUMMY_351 NETTRAN_DUMMY_352 BUF_X2 
XU28 IN4 n443 NETTRAN_DUMMY_353 NETTRAN_DUMMY_354 BUF_X2 
XU17 IN4 n442 NETTRAN_DUMMY_355 NETTRAN_DUMMY_356 BUF_X2 
XU12 IN4 n439 NETTRAN_DUMMY_357 NETTRAN_DUMMY_358 BUF_X2 
XU10 IN5 n435 NETTRAN_DUMMY_359 NETTRAN_DUMMY_360 BUF_X2 
XU2 n433 n434 NETTRAN_DUMMY_361 NETTRAN_DUMMY_362 INV_X1 
XU1 IN5 n433 NETTRAN_DUMMY_363 NETTRAN_DUMMY_364 BUF_X2 
XU66 n444 n14 n66 NETTRAN_DUMMY_365 NETTRAN_DUMMY_366 XOR2_X1 
XU65 n480 n458 n65 NETTRAN_DUMMY_367 NETTRAN_DUMMY_368 XOR2_X1 
XU64 n493 n1524 n64 NETTRAN_DUMMY_369 NETTRAN_DUMMY_370 XOR2_X1 
XU63 n493 n1536 n63 NETTRAN_DUMMY_371 NETTRAN_DUMMY_372 XOR2_X1 
XU62 n451 n1531 n62 NETTRAN_DUMMY_373 NETTRAN_DUMMY_374 XOR2_X1 
XU61 n488 n497 n61 NETTRAN_DUMMY_375 NETTRAN_DUMMY_376 XOR2_X1 
XU60 n468 n448 n60 NETTRAN_DUMMY_377 NETTRAN_DUMMY_378 XOR2_X1 
XU59 n1531 n1524 addr[5] n59 NETTRAN_DUMMY_379 NETTRAN_DUMMY_380 MUX2_X1 
XU57 n1531 addr[0] n448 n56 NETTRAN_DUMMY_381 NETTRAN_DUMMY_382 MUX2_X1 
XU54 n2 n1 addr[5] n53 NETTRAN_DUMMY_383 NETTRAN_DUMMY_384 MUX2_X1 
XU52 n1531 n1540 addr[5] n51 NETTRAN_DUMMY_385 NETTRAN_DUMMY_386 MUX2_X1 
XU51 n2 addr[0] addr[5] n50 NETTRAN_DUMMY_387 NETTRAN_DUMMY_388 MUX2_X1 
XU50 n6 n2 addr[5] n49 NETTRAN_DUMMY_389 NETTRAN_DUMMY_390 MUX2_X1 
XU48 n9 n1537 addr[5] n47 NETTRAN_DUMMY_391 NETTRAN_DUMMY_392 MUX2_X1 
XU45 n1540 n1524 addr[5] n44 NETTRAN_DUMMY_393 NETTRAN_DUMMY_394 MUX2_X1 
XU43 n1540 n501 n448 n42 NETTRAN_DUMMY_395 NETTRAN_DUMMY_396 MUX2_X1 
XU42 n1 n5 addr[5] n41 NETTRAN_DUMMY_397 NETTRAN_DUMMY_398 MUX2_X1 
XU41 n512 n1540 addr[5] n40 NETTRAN_DUMMY_399 NETTRAN_DUMMY_400 MUX2_X1 
XU40 addr[0] n1524 addr[5] n39 NETTRAN_DUMMY_401 NETTRAN_DUMMY_402 MUX2_X1 
XU38 n1540 n512 addr[5] n37 NETTRAN_DUMMY_403 NETTRAN_DUMMY_404 MUX2_X1 
XU36 n451 addr[1] n35 NETTRAN_DUMMY_405 NETTRAN_DUMMY_406 XOR2_X1 
XU35 n1531 n501 addr[5] n34 NETTRAN_DUMMY_407 NETTRAN_DUMMY_408 MUX2_X1 
XU34 addr[1] n1524 addr[5] n33 NETTRAN_DUMMY_409 NETTRAN_DUMMY_410 MUX2_X1 
XU33 n1524 n501 addr[5] n32 NETTRAN_DUMMY_411 NETTRAN_DUMMY_412 MUX2_X1 
XU32 n1531 addr[1] addr[5] n31 NETTRAN_DUMMY_413 NETTRAN_DUMMY_414 MUX2_X1 
XU31 n9 addr[0] addr[5] n30 NETTRAN_DUMMY_415 NETTRAN_DUMMY_416 MUX2_X1 
XU29 n2 addr[5] n28 NETTRAN_DUMMY_417 NETTRAN_DUMMY_418 XOR2_X1 
XU27 addr[0] n497 n448 n26 NETTRAN_DUMMY_419 NETTRAN_DUMMY_420 MUX2_X1 
XU26 n1537 n512 n448 n25 NETTRAN_DUMMY_421 NETTRAN_DUMMY_422 MUX2_X1 
XU25 n1537 addr[0] n448 n24 NETTRAN_DUMMY_423 NETTRAN_DUMMY_424 MUX2_X1 
XU24 n512 n2 n448 n23 NETTRAN_DUMMY_425 NETTRAN_DUMMY_426 MUX2_X1 
XU23 addr[0] n2 n448 n22 NETTRAN_DUMMY_427 NETTRAN_DUMMY_428 MUX2_X1 
XU21 n1527 addr[1] addr[5] n20 NETTRAN_DUMMY_429 NETTRAN_DUMMY_430 MUX2_X1 
XU19 n5 n501 n448 n18 NETTRAN_DUMMY_431 NETTRAN_DUMMY_432 MUX2_X1 
XU16 n501 addr[0] n9 NETTRAN_DUMMY_433 NETTRAN_DUMMY_434 XOR2_X1 
XU15 n1537 n1527 n448 n17 NETTRAN_DUMMY_435 NETTRAN_DUMMY_436 MUX2_X1 
Xc1_reg_0_ d[17] n63_G2B1I9 n2037 NETTRAN_DUMMY_437 NETTRAN_DUMMY_438 NETTRAN_DUMMY_439 DFF_X1 
Xc1_reg_1_ d[18] n63_G2B1I9 n2038 NETTRAN_DUMMY_440 NETTRAN_DUMMY_441 NETTRAN_DUMMY_442 DFF_X1 
Xc1_reg_2_ d[19] n63_G2B1I9 n2039 NETTRAN_DUMMY_443 NETTRAN_DUMMY_444 NETTRAN_DUMMY_445 DFF_X1 
Xc1_reg_3_ d[20] n63_G2B1I9 n2040 NETTRAN_DUMMY_446 NETTRAN_DUMMY_447 NETTRAN_DUMMY_448 DFF_X1 
Xc1_reg_4_ d[21] n63_G2B1I9 n2041 NETTRAN_DUMMY_449 NETTRAN_DUMMY_450 NETTRAN_DUMMY_451 DFF_X1 
Xc1_reg_5_ d[22] n63_G2B1I7 n2042 NETTRAN_DUMMY_452 NETTRAN_DUMMY_453 NETTRAN_DUMMY_454 DFF_X1 
Xc1_reg_6_ d[23] n63_G2B1I7 n2027 NETTRAN_DUMMY_455 NETTRAN_DUMMY_456 NETTRAN_DUMMY_457 DFF_X1 
Xc1_reg_7_ d[24] n63_G2B1I7 n2028 NETTRAN_DUMMY_458 NETTRAN_DUMMY_459 NETTRAN_DUMMY_460 DFF_X1 
Xc1_reg_8_ d[25] n63_G2B1I7 n2029 NETTRAN_DUMMY_461 NETTRAN_DUMMY_462 NETTRAN_DUMMY_463 DFF_X1 
Xc1_reg_9_ d[26] n63_G2B1I7 n2030 NETTRAN_DUMMY_464 NETTRAN_DUMMY_465 NETTRAN_DUMMY_466 DFF_X1 
Xc1_reg_10_ d[27] n63_G2B1I7 n2031 NETTRAN_DUMMY_467 NETTRAN_DUMMY_468 NETTRAN_DUMMY_469 DFF_X1 
Xc1_reg_11_ d[28] n63_G2B1I7 n2032 NETTRAN_DUMMY_470 NETTRAN_DUMMY_471 NETTRAN_DUMMY_472 DFF_X1 
Xc1_reg_12_ n457 clk_cts_1 n2033 NETTRAN_DUMMY_473 NETTRAN_DUMMY_474 NETTRAN_DUMMY_475 DFF_X1 
Xc1_reg_13_ d[30] clk_cts_1 n2034 NETTRAN_DUMMY_476 NETTRAN_DUMMY_477 NETTRAN_DUMMY_478 DFF_X1 
Xc1_reg_14_ n1548 clk_cts_0 n2019 NETTRAN_DUMMY_479 NETTRAN_DUMMY_480 NETTRAN_DUMMY_481 DFF_X1 
Xc1_reg_15_ n514 clk_cts_0 n2020 NETTRAN_DUMMY_482 NETTRAN_DUMMY_483 NETTRAN_DUMMY_484 DFF_X1 
Xc1_reg_16_ n2061 clk_cts_0 n2021 NETTRAN_DUMMY_485 NETTRAN_DUMMY_486 NETTRAN_DUMMY_487 DFF_X1 
Xc0_reg_0_ d[35] n63_G2B1I6 n2051 NETTRAN_DUMMY_488 NETTRAN_DUMMY_489 NETTRAN_DUMMY_490 DFF_X1 
Xc0_reg_1_ d[36] n63_G2B1I6 n2052 NETTRAN_DUMMY_491 NETTRAN_DUMMY_492 NETTRAN_DUMMY_493 DFF_X1 
Xc0_reg_2_ d[37] n63_G2B1I6 n2053 NETTRAN_DUMMY_494 NETTRAN_DUMMY_495 NETTRAN_DUMMY_496 DFF_X1 
Xc0_reg_3_ d[38] n63_G2B1I6 n2054 NETTRAN_DUMMY_497 NETTRAN_DUMMY_498 NETTRAN_DUMMY_499 DFF_X1 
Xc0_reg_4_ d[39] n63_G2B1I5 n2055 NETTRAN_DUMMY_500 NETTRAN_DUMMY_501 NETTRAN_DUMMY_502 DFF_X1 
Xc0_reg_5_ d[40] n63_G2B1I5 n2056 NETTRAN_DUMMY_503 NETTRAN_DUMMY_504 NETTRAN_DUMMY_505 DFF_X1 
Xc0_reg_6_ d[41] n63_G2B1I5 n2057 NETTRAN_DUMMY_506 NETTRAN_DUMMY_507 NETTRAN_DUMMY_508 DFF_X1 
Xc0_reg_7_ d[42] n63_G2B1I6 n2058 NETTRAN_DUMMY_509 NETTRAN_DUMMY_510 NETTRAN_DUMMY_511 DFF_X1 
Xc0_reg_8_ d[43] n63_G2B1I5 n2043 NETTRAN_DUMMY_512 NETTRAN_DUMMY_513 NETTRAN_DUMMY_514 DFF_X1 
Xc0_reg_9_ n506 clk_cts_1 n2044 NETTRAN_DUMMY_515 NETTRAN_DUMMY_516 NETTRAN_DUMMY_517 DFF_X1 
Xc0_reg_10_ n504 clk_cts_0 n2045 NETTRAN_DUMMY_518 NETTRAN_DUMMY_519 NETTRAN_DUMMY_520 DFF_X1 
Xc0_reg_11_ n498 n63_G2B1I9 n2046 NETTRAN_DUMMY_521 NETTRAN_DUMMY_522 NETTRAN_DUMMY_523 DFF_X1 
Xc0_reg_12_ n496 n63_G2B1I9 n2047 NETTRAN_DUMMY_524 NETTRAN_DUMMY_525 NETTRAN_DUMMY_526 DFF_X1 
Xc0_reg_13_ n494 n63_G2B1I9 n2048 NETTRAN_DUMMY_527 NETTRAN_DUMMY_528 NETTRAN_DUMMY_529 DFF_X1 
Xc0_reg_14_ n490 n63_G2B1I6 n2049 NETTRAN_DUMMY_530 NETTRAN_DUMMY_531 NETTRAN_DUMMY_532 DFF_X1 
Xc0_reg_15_ n2060 n63_G2B1I1 n2050 NETTRAN_DUMMY_533 NETTRAN_DUMMY_534 NETTRAN_DUMMY_535 DFF_X1 
Xc0_reg_16_ N4680 n63_G2B1I6 n2035 NETTRAN_DUMMY_536 NETTRAN_DUMMY_537 NETTRAN_DUMMY_538 DFF_X1 
Xc0_reg_17_ N4640 n63_G2B1I1 n2036 NETTRAN_DUMMY_539 NETTRAN_DUMMY_540 NETTRAN_DUMMY_541 DFF_X1 
Xc2_reg_0_ d[0] n63_G2B1I4 n2023 NETTRAN_DUMMY_542 NETTRAN_DUMMY_543 NETTRAN_DUMMY_544 DFF_X1 
Xc2_reg_1_ d[1] clk_cts_0 n2024 NETTRAN_DUMMY_545 NETTRAN_DUMMY_546 NETTRAN_DUMMY_547 DFF_X1 
Xc2_reg_2_ d[2] n63_G2B1I1 n2025 NETTRAN_DUMMY_548 NETTRAN_DUMMY_549 NETTRAN_DUMMY_550 DFF_X1 
Xc2_reg_3_ d[3] n63_G2B1I9 n2026 NETTRAN_DUMMY_551 NETTRAN_DUMMY_552 NETTRAN_DUMMY_553 DFF_X1 
Xc2_reg_4_ d[4] n63_G2B1I3 n2011 NETTRAN_DUMMY_554 NETTRAN_DUMMY_555 NETTRAN_DUMMY_556 DFF_X1 
Xc2_reg_5_ n478 n63_G2B1I3 n2012 NETTRAN_DUMMY_557 NETTRAN_DUMMY_558 NETTRAN_DUMMY_559 DFF_X1 
Xc2_reg_6_ n474 n63_G2B1I3 n2013 NETTRAN_DUMMY_560 NETTRAN_DUMMY_561 NETTRAN_DUMMY_562 DFF_X1 
Xc2_reg_7_ d[7] n63_G2B1I1 n2014 NETTRAN_DUMMY_563 NETTRAN_DUMMY_564 NETTRAN_DUMMY_565 DFF_X1 
Xc2_reg_8_ n470 n63_G2B1I3 n2015 NETTRAN_DUMMY_566 NETTRAN_DUMMY_567 NETTRAN_DUMMY_568 DFF_X1 
Xc2_reg_9_ n467 n63_G2B1I3 n2016 NETTRAN_DUMMY_569 NETTRAN_DUMMY_570 NETTRAN_DUMMY_571 DFF_X1 
Xc2_reg_10_ d[10] n63_G2B1I4 n2017 NETTRAN_DUMMY_572 NETTRAN_DUMMY_573 NETTRAN_DUMMY_574 DFF_X1 
Xc2_reg_11_ d[11] n63_G2B1I4 n2018 NETTRAN_DUMMY_575 NETTRAN_DUMMY_576 NETTRAN_DUMMY_577 DFF_X1 
Xc2_reg_12_ d[12] n63_G2B1I4 n2006 NETTRAN_DUMMY_578 NETTRAN_DUMMY_579 NETTRAN_DUMMY_580 DFF_X1 
Xc2_reg_13_ d[13] n63_G2B1I4 n2007 NETTRAN_DUMMY_581 NETTRAN_DUMMY_582 NETTRAN_DUMMY_583 DFF_X1 
Xc2_reg_14_ d[14] n63_G2B1I4 n2008 NETTRAN_DUMMY_584 NETTRAN_DUMMY_585 NETTRAN_DUMMY_586 DFF_X1 
Xc2_reg_15_ n459 n63_G2B1I4 n2009 NETTRAN_DUMMY_587 NETTRAN_DUMMY_588 NETTRAN_DUMMY_589 DFF_X1 
Xc2_reg_16_ N19520 n63_G2B1I4 n2010 NETTRAN_DUMMY_590 NETTRAN_DUMMY_591 NETTRAN_DUMMY_592 DFF_X1 
XU162 n160 n151 addr[7] n161 NETTRAN_DUMMY_593 NETTRAN_DUMMY_594 MUX2_X1 
XU161 n159 n155 addr[4] n160 NETTRAN_DUMMY_595 NETTRAN_DUMMY_596 MUX2_X1 
XU160 n158 n156 addr[3] n159 NETTRAN_DUMMY_597 NETTRAN_DUMMY_598 MUX2_X1 
XU159 n157 n1630 addr[2] n158 NETTRAN_DUMMY_599 NETTRAN_DUMMY_600 MUX2_X1 
XU158 n1 addr[1] addr[5] n157 NETTRAN_DUMMY_601 NETTRAN_DUMMY_602 MUX2_X1 
XU157 n1631 n1632 addr[2] n156 NETTRAN_DUMMY_603 NETTRAN_DUMMY_604 MUX2_X1 
XU156 n154 n152 addr[3] n155 NETTRAN_DUMMY_605 NETTRAN_DUMMY_606 MUX2_X1 
XU155 n153 n62 addr[2] n154 NETTRAN_DUMMY_607 NETTRAN_DUMMY_608 MUX2_X1 
XU154 n2 addr[1] addr[5] n153 NETTRAN_DUMMY_609 NETTRAN_DUMMY_610 MUX2_X1 
XU153 n1648 n1628 addr[2] n152 NETTRAN_DUMMY_611 NETTRAN_DUMMY_612 MUX2_X1 
XU152 n150 n147 addr[4] n151 NETTRAN_DUMMY_613 NETTRAN_DUMMY_614 MUX2_X1 
XU151 n149 n148 n484 n150 NETTRAN_DUMMY_615 NETTRAN_DUMMY_616 MUX2_X1 
XU150 n11 n1597 addr[2] n149 NETTRAN_DUMMY_617 NETTRAN_DUMMY_618 MUX2_X1 
XU149 n32 n5 addr[2] n148 NETTRAN_DUMMY_619 NETTRAN_DUMMY_620 MUX2_X1 
XU148 n146 n145 n484 n147 NETTRAN_DUMMY_621 NETTRAN_DUMMY_622 MUX2_X1 
XU146 addr[1] n1596 IN0 n145 NETTRAN_DUMMY_623 NETTRAN_DUMMY_624 MUX2_X1 
XU145 n143 n138 addr[7] n144 NETTRAN_DUMMY_625 NETTRAN_DUMMY_626 MUX2_X1 
XU144 n142 n140 n458 n143 NETTRAN_DUMMY_627 NETTRAN_DUMMY_628 MUX2_X1 
XU143 n141 n64 n484 n142 NETTRAN_DUMMY_629 NETTRAN_DUMMY_630 MUX2_X1 
XU142 n1633 n1634 IN0 n141 NETTRAN_DUMMY_631 NETTRAN_DUMMY_632 MUX2_X1 
XU141 n139 n63 n484 n140 NETTRAN_DUMMY_633 NETTRAN_DUMMY_634 MUX2_X1 
XU140 n5 n1596 IN0 n139 NETTRAN_DUMMY_635 NETTRAN_DUMMY_636 MUX2_X1 
XU139 n137 n135 n458 n138 NETTRAN_DUMMY_637 NETTRAN_DUMMY_638 MUX2_X1 
XU138 n449 n136 n429 n137 NETTRAN_DUMMY_639 NETTRAN_DUMMY_640 MUX2_X1 
XU137 n12 n411 n480 n136 NETTRAN_DUMMY_641 NETTRAN_DUMMY_642 MUX2_X1 
XU136 n134 n1598 n484 n135 NETTRAN_DUMMY_643 NETTRAN_DUMMY_644 MUX2_X1 
XU135 n1655 n430 IN0 n134 NETTRAN_DUMMY_645 NETTRAN_DUMMY_646 MUX2_X1 
XU134 n133 n116 addr[6] d[45] NETTRAN_DUMMY_647 NETTRAN_DUMMY_648 MUX2_X1 
XU133 n132 n123 addr[7] n133 NETTRAN_DUMMY_649 NETTRAN_DUMMY_650 MUX2_X1 
XU132 n131 n126 addr[4] n132 NETTRAN_DUMMY_651 NETTRAN_DUMMY_652 MUX2_X1 
XU131 n128 n129 addr[2] n131 NETTRAN_DUMMY_653 NETTRAN_DUMMY_654 MUX2_X1 
XU129 n1624 n127 addr[3] n128 NETTRAN_DUMMY_655 NETTRAN_DUMMY_656 MUX2_X1 
XU128 addr[1] n9 addr[5] n127 NETTRAN_DUMMY_657 NETTRAN_DUMMY_658 MUX2_X1 
XU127 n125 n124 IN0 n126 NETTRAN_DUMMY_659 NETTRAN_DUMMY_660 MUX2_X1 
XU126 n1645 n1651 n487 n125 NETTRAN_DUMMY_661 NETTRAN_DUMMY_662 MUX2_X1 
XU125 addr[0] n22 n487 n124 NETTRAN_DUMMY_663 NETTRAN_DUMMY_664 MUX2_X1 
XU124 n122 n119 addr[4] n123 NETTRAN_DUMMY_665 NETTRAN_DUMMY_666 MUX2_X1 
XU123 n121 n120 addr[2] n122 NETTRAN_DUMMY_667 NETTRAN_DUMMY_668 MUX2_X1 
XU122 n1625 n1626 addr[3] n121 NETTRAN_DUMMY_669 NETTRAN_DUMMY_670 MUX2_X1 
XU121 n33 n8 addr[3] n120 NETTRAN_DUMMY_671 NETTRAN_DUMMY_672 MUX2_X1 
XU120 n61 n118 IN0 n119 NETTRAN_DUMMY_673 NETTRAN_DUMMY_674 MUX2_X1 
XU119 n9 n117 n484 n118 NETTRAN_DUMMY_675 NETTRAN_DUMMY_676 MUX2_X1 
XU118 n5 n6 n448 n117 NETTRAN_DUMMY_677 NETTRAN_DUMMY_678 MUX2_X1 
XU117 n115 n108 addr[7] n116 NETTRAN_DUMMY_679 NETTRAN_DUMMY_680 MUX2_X1 
XU116 n114 n111 addr[4] n115 NETTRAN_DUMMY_681 NETTRAN_DUMMY_682 MUX2_X1 
XU115 n113 n112 addr[2] n114 NETTRAN_DUMMY_683 NETTRAN_DUMMY_684 MUX2_X1 
XU114 n1628 n27 addr[3] n113 NETTRAN_DUMMY_685 NETTRAN_DUMMY_686 MUX2_X1 
XU113 n1627 n1531 addr[3] n112 NETTRAN_DUMMY_687 NETTRAN_DUMMY_688 MUX2_X1 
XU112 n110 n109 addr[2] n111 NETTRAN_DUMMY_689 NETTRAN_DUMMY_690 MUX2_X1 
XU111 n1531 n1595 addr[3] n110 NETTRAN_DUMMY_691 NETTRAN_DUMMY_692 MUX2_X1 
XU110 n34 n33 addr[3] n109 NETTRAN_DUMMY_693 NETTRAN_DUMMY_694 MUX2_X1 
XU109 n107 n103 addr[4] n108 NETTRAN_DUMMY_695 NETTRAN_DUMMY_696 MUX2_X1 
XU108 n106 n104 addr[2] n107 NETTRAN_DUMMY_697 NETTRAN_DUMMY_698 MUX2_X1 
XU107 n105 n8 addr[3] n106 NETTRAN_DUMMY_699 NETTRAN_DUMMY_700 MUX2_X1 
XU105 n33 n32 addr[3] n104 NETTRAN_DUMMY_701 NETTRAN_DUMMY_702 MUX2_X1 
XU104 n102 n101 addr[2] n103 NETTRAN_DUMMY_703 NETTRAN_DUMMY_704 MUX2_X1 
XU103 n1654 n1596 n484 n102 NETTRAN_DUMMY_705 NETTRAN_DUMMY_706 MUX2_X1 
XU102 n1629 n1597 n484 n101 NETTRAN_DUMMY_707 NETTRAN_DUMMY_708 MUX2_X1 
XU101 n100 n83 n445 d[44] NETTRAN_DUMMY_709 NETTRAN_DUMMY_710 MUX2_X1 
XU100 n99 n91 n433 n100 NETTRAN_DUMMY_711 NETTRAN_DUMMY_712 MUX2_X1 
XU99 n98 n94 IN0 n99 NETTRAN_DUMMY_713 NETTRAN_DUMMY_714 MUX2_X1 
XU98 n97 n95 n487 n98 NETTRAN_DUMMY_715 NETTRAN_DUMMY_716 MUX2_X1 
XU97 n1609 n96 n460 n97 NETTRAN_DUMMY_717 NETTRAN_DUMMY_718 MUX2_X1 
XU96 n497 n1531 n448 n96 NETTRAN_DUMMY_719 NETTRAN_DUMMY_720 MUX2_X1 
XU95 n1653 n3 n460 n95 NETTRAN_DUMMY_721 NETTRAN_DUMMY_722 MUX2_X1 
XU94 n93 n92 n487 n94 NETTRAN_DUMMY_723 NETTRAN_DUMMY_724 MUX2_X1 
XU93 n1614 n1613 n460 n93 NETTRAN_DUMMY_725 NETTRAN_DUMMY_726 MUX2_X1 
XU92 n1616 n1617 n460 n92 NETTRAN_DUMMY_727 NETTRAN_DUMMY_728 MUX2_X1 
XU91 n90 n86 IN0 n91 NETTRAN_DUMMY_729 NETTRAN_DUMMY_730 MUX2_X1 
XU90 n89 n88 n487 n90 NETTRAN_DUMMY_731 NETTRAN_DUMMY_732 MUX2_X1 
XU89 n22 n23 n460 n89 NETTRAN_DUMMY_733 NETTRAN_DUMMY_734 MUX2_X1 
XU88 n87 n2 n60 n88 NETTRAN_DUMMY_735 NETTRAN_DUMMY_736 MUX2_X1 
XU87 n1527 n512 n468 n87 NETTRAN_DUMMY_737 NETTRAN_DUMMY_738 MUX2_X1 
XU86 n85 n84 n487 n86 NETTRAN_DUMMY_739 NETTRAN_DUMMY_740 MUX2_X1 
XU85 n1618 addr[0] n460 n85 NETTRAN_DUMMY_741 NETTRAN_DUMMY_742 MUX2_X1 
XU84 n1619 n1652 n460 n84 NETTRAN_DUMMY_743 NETTRAN_DUMMY_744 MUX2_X1 
XU83 n82 n75 n433 n83 NETTRAN_DUMMY_745 NETTRAN_DUMMY_746 MUX2_X1 
XU82 n81 n78 IN0 n82 NETTRAN_DUMMY_747 NETTRAN_DUMMY_748 MUX2_X1 
XU81 n80 n79 n487 n81 NETTRAN_DUMMY_749 NETTRAN_DUMMY_750 MUX2_X1 
XU80 n1620 n1621 n460 n80 NETTRAN_DUMMY_751 NETTRAN_DUMMY_752 MUX2_X1 
XU79 n24 n512 n460 n79 NETTRAN_DUMMY_753 NETTRAN_DUMMY_754 MUX2_X1 
XU78 n77 n76 n487 n78 NETTRAN_DUMMY_755 NETTRAN_DUMMY_756 MUX2_X1 
XU77 n1622 n1620 n460 n77 NETTRAN_DUMMY_757 NETTRAN_DUMMY_758 MUX2_X1 
XU76 addr[0] n1618 n460 n76 NETTRAN_DUMMY_759 NETTRAN_DUMMY_760 MUX2_X1 
XU75 n74 n71 IN0 n75 NETTRAN_DUMMY_761 NETTRAN_DUMMY_762 MUX2_X1 
XU74 n73 n72 n487 n74 NETTRAN_DUMMY_763 NETTRAN_DUMMY_764 MUX2_X1 
XU73 n1652 n1607 n460 n73 NETTRAN_DUMMY_765 NETTRAN_DUMMY_766 MUX2_X1 
XU72 n1651 n1602 n468 n72 NETTRAN_DUMMY_767 NETTRAN_DUMMY_768 MUX2_X1 
XU71 n1604 n70 n487 n71 NETTRAN_DUMMY_769 NETTRAN_DUMMY_770 MUX2_X1 
XU70 n1645 n1594 n460 n70 NETTRAN_DUMMY_771 NETTRAN_DUMMY_772 MUX2_X1 
XU69 n449 n1 n69 NETTRAN_DUMMY_773 NETTRAN_DUMMY_774 XOR2_X1 
XU68 n448 n433 n68 NETTRAN_DUMMY_775 NETTRAN_DUMMY_776 XOR2_X1 
XU67 n480 n433 n67 NETTRAN_DUMMY_777 NETTRAN_DUMMY_778 XOR2_X1 
XU273 n27 n271 n433 n272 NETTRAN_DUMMY_779 NETTRAN_DUMMY_780 MUX2_X1 
XU272 n501 n1537 n448 n271 NETTRAN_DUMMY_781 NETTRAN_DUMMY_782 MUX2_X1 
XU271 n269 n1524 n68 n270 NETTRAN_DUMMY_783 NETTRAN_DUMMY_784 MUX2_X1 
XU270 n5 n1537 n433 n269 NETTRAN_DUMMY_785 NETTRAN_DUMMY_786 MUX2_X1 
XU269 n267 n266 n487 n268 NETTRAN_DUMMY_787 NETTRAN_DUMMY_788 MUX2_X1 
XU267 n1658 n26 addr[7] n266 NETTRAN_DUMMY_789 NETTRAN_DUMMY_790 MUX2_X1 
XU266 n264 n260 addr[2] n265 NETTRAN_DUMMY_791 NETTRAN_DUMMY_792 MUX2_X1 
XU265 n263 n262 n487 n264 NETTRAN_DUMMY_793 NETTRAN_DUMMY_794 MUX2_X1 
XU264 n47 n1 addr[7] n263 NETTRAN_DUMMY_795 NETTRAN_DUMMY_796 MUX2_X1 
XU263 n58 n261 addr[7] n262 NETTRAN_DUMMY_797 NETTRAN_DUMMY_798 MUX2_X1 
XU260 n258 n259 n487 n260 NETTRAN_DUMMY_799 NETTRAN_DUMMY_800 MUX2_X1 
XU258 n1656 n1657 addr[7] n258 NETTRAN_DUMMY_801 NETTRAN_DUMMY_802 MUX2_X1 
XU257 n256 n250 n460 n257 NETTRAN_DUMMY_803 NETTRAN_DUMMY_804 MUX2_X1 
XU256 n255 n253 n492 n256 NETTRAN_DUMMY_805 NETTRAN_DUMMY_806 MUX2_X1 
XU255 n254 n1655 n67 n255 NETTRAN_DUMMY_807 NETTRAN_DUMMY_808 MUX2_X1 
XU254 n43 n1640 n484 n254 NETTRAN_DUMMY_809 NETTRAN_DUMMY_810 MUX2_X1 
XU253 n252 n251 n487 n253 NETTRAN_DUMMY_811 NETTRAN_DUMMY_812 MUX2_X1 
XU251 n1615 n1536 n433 n251 NETTRAN_DUMMY_813 NETTRAN_DUMMY_814 MUX2_X1 
XU250 n249 n245 IN0 n250 NETTRAN_DUMMY_815 NETTRAN_DUMMY_816 MUX2_X1 
XU249 n247 n246 n484 n249 NETTRAN_DUMMY_817 NETTRAN_DUMMY_818 MUX2_X1 
XU247 n1650 n1597 addr[7] n246 NETTRAN_DUMMY_819 NETTRAN_DUMMY_820 MUX2_X1 
XU246 n244 n242 n484 n245 NETTRAN_DUMMY_821 NETTRAN_DUMMY_822 MUX2_X1 
XU245 n243 n1605 addr[7] n244 NETTRAN_DUMMY_823 NETTRAN_DUMMY_824 MUX2_X1 
XU244 n501 n1524 n455 n243 NETTRAN_DUMMY_825 NETTRAN_DUMMY_826 MUX2_X1 
XU243 n1606 n1591 addr[7] n242 NETTRAN_DUMMY_827 NETTRAN_DUMMY_828 MUX2_X1 
XU242 n241 n225 addr[6] d[4] NETTRAN_DUMMY_829 NETTRAN_DUMMY_830 MUX2_X1 
XU241 n240 n232 addr[7] n241 NETTRAN_DUMMY_831 NETTRAN_DUMMY_832 MUX2_X1 
XU240 n239 n234 addr[4] n240 NETTRAN_DUMMY_833 NETTRAN_DUMMY_834 MUX2_X1 
XU239 n238 n237 addr[2] n239 NETTRAN_DUMMY_835 NETTRAN_DUMMY_836 MUX2_X1 
XU238 n1631 n1637 addr[3] n238 NETTRAN_DUMMY_837 NETTRAN_DUMMY_838 MUX2_X1 
XU237 n236 n235 addr[3] n237 NETTRAN_DUMMY_839 NETTRAN_DUMMY_840 MUX2_X1 
XU236 n2 n6 addr[5] n236 NETTRAN_DUMMY_841 NETTRAN_DUMMY_842 MUX2_X1 
XU235 n1527 n1524 addr[5] n235 NETTRAN_DUMMY_843 NETTRAN_DUMMY_844 MUX2_X1 
XU234 n233 n1597 addr[2] n234 NETTRAN_DUMMY_845 NETTRAN_DUMMY_846 MUX2_X1 
XU233 n1611 n512 n487 n233 NETTRAN_DUMMY_847 NETTRAN_DUMMY_848 MUX2_X1 
XU232 n231 n228 addr[4] n232 NETTRAN_DUMMY_849 NETTRAN_DUMMY_850 MUX2_X1 
XU231 n230 n229 addr[2] n231 NETTRAN_DUMMY_851 NETTRAN_DUMMY_852 MUX2_X1 
XU230 n37 n15 addr[3] n230 NETTRAN_DUMMY_853 NETTRAN_DUMMY_854 MUX2_X1 
XU229 n26 n39 addr[3] n229 NETTRAN_DUMMY_855 NETTRAN_DUMMY_856 MUX2_X1 
XU228 n227 n226 addr[2] n228 NETTRAN_DUMMY_857 NETTRAN_DUMMY_858 MUX2_X1 
XU227 n411 n1638 n487 n227 NETTRAN_DUMMY_859 NETTRAN_DUMMY_860 MUX2_X1 
XU226 n30 n1639 addr[3] n226 NETTRAN_DUMMY_861 NETTRAN_DUMMY_862 MUX2_X1 
XU225 n224 n216 addr[7] n225 NETTRAN_DUMMY_863 NETTRAN_DUMMY_864 MUX2_X1 
XU224 n222 n219 addr[4] n224 NETTRAN_DUMMY_865 NETTRAN_DUMMY_866 MUX2_X1 
XU222 n221 n1611 addr[2] n220 NETTRAN_DUMMY_867 NETTRAN_DUMMY_868 MUX2_X1 
XU221 n218 n217 addr[2] n219 NETTRAN_DUMMY_869 NETTRAN_DUMMY_870 MUX2_X1 
XU220 n7 n1640 addr[3] n218 NETTRAN_DUMMY_871 NETTRAN_DUMMY_872 MUX2_X1 
XU219 n6 n1599 n484 n217 NETTRAN_DUMMY_873 NETTRAN_DUMMY_874 MUX2_X1 
XU218 n215 n212 addr[4] n216 NETTRAN_DUMMY_875 NETTRAN_DUMMY_876 MUX2_X1 
XU217 n214 n213 addr[2] n215 NETTRAN_DUMMY_877 NETTRAN_DUMMY_878 MUX2_X1 
XU216 n427 n1591 n484 n214 NETTRAN_DUMMY_879 NETTRAN_DUMMY_880 MUX2_X1 
XU215 n105 n1594 n484 n213 NETTRAN_DUMMY_881 NETTRAN_DUMMY_882 MUX2_X1 
XU214 n211 n210 n492 n212 NETTRAN_DUMMY_883 NETTRAN_DUMMY_884 MUX2_X1 
XU212 n1605 n449 n484 n210 NETTRAN_DUMMY_885 NETTRAN_DUMMY_886 MUX2_X1 
XU211 n209 n196 addr[7] d[48] NETTRAN_DUMMY_887 NETTRAN_DUMMY_888 MUX2_X1 
XU210 n208 n202 n458 n209 NETTRAN_DUMMY_889 NETTRAN_DUMMY_890 MUX2_X1 
XU209 n206 n207 IN0 n208 NETTRAN_DUMMY_891 NETTRAN_DUMMY_892 MUX2_X1 
XU207 n205 n203 n445 n206 NETTRAN_DUMMY_893 NETTRAN_DUMMY_894 MUX2_X1 
XU204 n199 n200 IN0 n202 NETTRAN_DUMMY_895 NETTRAN_DUMMY_896 MUX2_X1 
XU202 n197 n198 n445 n199 NETTRAN_DUMMY_897 NETTRAN_DUMMY_898 MUX2_X1 
XU200 n12 n427 n480 n197 NETTRAN_DUMMY_899 NETTRAN_DUMMY_900 MUX2_X1 
XU199 n195 n191 n458 n196 NETTRAN_DUMMY_901 NETTRAN_DUMMY_902 MUX2_X1 
XU198 n66 n194 IN0 n195 NETTRAN_DUMMY_903 NETTRAN_DUMMY_904 MUX2_X1 
XU197 n193 n192 n445 n194 NETTRAN_DUMMY_905 NETTRAN_DUMMY_906 MUX2_X1 
XU195 n12 n455 n480 n192 NETTRAN_DUMMY_907 NETTRAN_DUMMY_908 MUX2_X1 
XU194 n190 n187 IN0 n191 NETTRAN_DUMMY_909 NETTRAN_DUMMY_910 MUX2_X1 
XU193 n189 n188 n445 n190 NETTRAN_DUMMY_911 NETTRAN_DUMMY_912 MUX2_X1 
XU190 n14 n186 n445 n187 NETTRAN_DUMMY_913 NETTRAN_DUMMY_914 MUX2_X1 
XU189 n1636 n1536 n484 n186 NETTRAN_DUMMY_915 NETTRAN_DUMMY_916 MUX2_X1 
XU188 n185 n171 n445 d[47] NETTRAN_DUMMY_917 NETTRAN_DUMMY_918 MUX2_X1 
XU187 n184 n177 addr[7] n185 NETTRAN_DUMMY_919 NETTRAN_DUMMY_920 MUX2_X1 
XU186 n183 n180 addr[4] n184 NETTRAN_DUMMY_921 NETTRAN_DUMMY_922 MUX2_X1 
XU185 n182 n181 n484 n183 NETTRAN_DUMMY_923 NETTRAN_DUMMY_924 MUX2_X1 
XU184 n31 n33 addr[2] n182 NETTRAN_DUMMY_925 NETTRAN_DUMMY_926 MUX2_X1 
XU183 n13 n1536 IN0 n181 NETTRAN_DUMMY_927 NETTRAN_DUMMY_928 MUX2_X1 
XU182 n179 n178 n484 n180 NETTRAN_DUMMY_929 NETTRAN_DUMMY_930 MUX2_X1 
XU181 n1595 n1635 addr[2] n179 NETTRAN_DUMMY_931 NETTRAN_DUMMY_932 MUX2_X1 
XU180 n1591 n1656 addr[2] n178 NETTRAN_DUMMY_933 NETTRAN_DUMMY_934 MUX2_X1 
XU179 n176 n173 n458 n177 NETTRAN_DUMMY_935 NETTRAN_DUMMY_936 MUX2_X1 
XU178 n175 n174 n480 n176 NETTRAN_DUMMY_937 NETTRAN_DUMMY_938 MUX2_X1 
XU177 n449 n12 IN0 n175 NETTRAN_DUMMY_939 NETTRAN_DUMMY_940 MUX2_X1 
XU176 n455 n411 IN0 n174 NETTRAN_DUMMY_941 NETTRAN_DUMMY_942 MUX2_X1 
XU175 n449 n172 n484 n173 NETTRAN_DUMMY_943 NETTRAN_DUMMY_944 MUX2_X1 
XU174 n1595 n455 IN0 n172 NETTRAN_DUMMY_945 NETTRAN_DUMMY_946 MUX2_X1 
XU173 n170 n165 addr[7] n171 NETTRAN_DUMMY_947 NETTRAN_DUMMY_948 MUX2_X1 
XU172 n169 n167 n458 n170 NETTRAN_DUMMY_949 NETTRAN_DUMMY_950 MUX2_X1 
XU171 n168 n45 n480 n169 NETTRAN_DUMMY_951 NETTRAN_DUMMY_952 MUX2_X1 
XU169 n1851 n166 n480 n167 NETTRAN_DUMMY_953 NETTRAN_DUMMY_954 MUX2_X1 
XU167 n1598 n164 n65 n165 NETTRAN_DUMMY_955 NETTRAN_DUMMY_956 MUX2_X1 
XU166 n163 n162 n458 n164 NETTRAN_DUMMY_957 NETTRAN_DUMMY_958 MUX2_X1 
XU165 n1634 n455 n492 n163 NETTRAN_DUMMY_959 NETTRAN_DUMMY_960 MUX2_X1 
XU164 n38 n19 n492 n162 NETTRAN_DUMMY_961 NETTRAN_DUMMY_962 MUX2_X1 
XU163 n161 n144 addr[6] d[46] NETTRAN_DUMMY_963 NETTRAN_DUMMY_964 MUX2_X1 
XU376 n374 n366 n460 n375 NETTRAN_DUMMY_965 NETTRAN_DUMMY_966 MUX2_X1 
XU375 n373 n369 addr[2] n374 NETTRAN_DUMMY_967 NETTRAN_DUMMY_968 MUX2_X1 
XU374 n372 n370 n487 n373 NETTRAN_DUMMY_969 NETTRAN_DUMMY_970 MUX2_X1 
XU373 n16 n371 addr[7] n372 NETTRAN_DUMMY_971 NETTRAN_DUMMY_972 MUX2_X1 
XU372 addr[0] n1540 addr[5] n371 NETTRAN_DUMMY_973 NETTRAN_DUMMY_974 MUX2_X1 
XU371 addr[1] n1658 addr[7] n370 NETTRAN_DUMMY_975 NETTRAN_DUMMY_976 MUX2_X1 
XU370 n368 n367 n487 n369 NETTRAN_DUMMY_977 NETTRAN_DUMMY_978 MUX2_X1 
XU369 n9 n46 addr[7] n368 NETTRAN_DUMMY_979 NETTRAN_DUMMY_980 MUX2_X1 
XU368 n1617 n19 addr[7] n367 NETTRAN_DUMMY_981 NETTRAN_DUMMY_982 MUX2_X1 
XU367 n365 n361 addr[2] n366 NETTRAN_DUMMY_983 NETTRAN_DUMMY_984 MUX2_X1 
XU366 n364 n362 n487 n365 NETTRAN_DUMMY_985 NETTRAN_DUMMY_986 MUX2_X1 
XU365 n363 n12 addr[7] n364 NETTRAN_DUMMY_987 NETTRAN_DUMMY_988 MUX2_X1 
XU364 n6 n1 n448 n363 NETTRAN_DUMMY_989 NETTRAN_DUMMY_990 MUX2_X1 
XU363 n3 n1622 addr[7] n362 NETTRAN_DUMMY_991 NETTRAN_DUMMY_992 MUX2_X1 
XU362 n360 n359 n487 n361 NETTRAN_DUMMY_993 NETTRAN_DUMMY_994 MUX2_X1 
XU361 n41 n20 addr[7] n360 NETTRAN_DUMMY_995 NETTRAN_DUMMY_996 MUX2_X1 
XU360 n36 n358 addr[7] n359 NETTRAN_DUMMY_997 NETTRAN_DUMMY_998 MUX2_X1 
XU358 n356 n348 n460 n357 NETTRAN_DUMMY_999 NETTRAN_DUMMY_1000 MUX2_X1 
XU357 n355 n352 IN0 n356 NETTRAN_DUMMY_1001 NETTRAN_DUMMY_1002 MUX2_X1 
XU356 n353 n354 n487 n355 NETTRAN_DUMMY_1003 NETTRAN_DUMMY_1004 MUX2_X1 
XU354 n1638 n1607 addr[7] n353 NETTRAN_DUMMY_1005 NETTRAN_DUMMY_1006 MUX2_X1 
XU353 n350 n351 n487 n352 NETTRAN_DUMMY_1007 NETTRAN_DUMMY_1008 MUX2_X1 
XU351 n52 n349 addr[7] n350 NETTRAN_DUMMY_1009 NETTRAN_DUMMY_1010 MUX2_X1 
XU350 n5 n9 n448 n349 NETTRAN_DUMMY_1011 NETTRAN_DUMMY_1012 MUX2_X1 
XU349 n345 n346 IN0 n348 NETTRAN_DUMMY_1013 NETTRAN_DUMMY_1014 MUX2_X1 
XU347 n344 n343 n484 n345 NETTRAN_DUMMY_1015 NETTRAN_DUMMY_1016 MUX2_X1 
XU346 n1605 n1599 addr[7] n344 NETTRAN_DUMMY_1017 NETTRAN_DUMMY_1018 MUX2_X1 
XU345 n56 n342 addr[7] n343 NETTRAN_DUMMY_1019 NETTRAN_DUMMY_1020 MUX2_X1 
XU343 n430 n69 n480 n341 NETTRAN_DUMMY_1021 NETTRAN_DUMMY_1022 MUX2_X1 
XU342 n340 n324 addr[6] d[7] NETTRAN_DUMMY_1023 NETTRAN_DUMMY_1024 MUX2_X1 
XU341 n339 n332 addr[7] n340 NETTRAN_DUMMY_1025 NETTRAN_DUMMY_1026 MUX2_X1 
XU340 n338 n335 addr[4] n339 NETTRAN_DUMMY_1027 NETTRAN_DUMMY_1028 MUX2_X1 
XU339 n337 n336 addr[2] n338 NETTRAN_DUMMY_1029 NETTRAN_DUMMY_1030 MUX2_X1 
XU338 n1603 n31 n484 n337 NETTRAN_DUMMY_1031 NETTRAN_DUMMY_1032 MUX2_X1 
XU337 n1599 n5 n484 n336 NETTRAN_DUMMY_1033 NETTRAN_DUMMY_1034 MUX2_X1 
XU336 n334 n333 addr[2] n335 NETTRAN_DUMMY_1035 NETTRAN_DUMMY_1036 MUX2_X1 
XU335 n56 n1608 n484 n334 NETTRAN_DUMMY_1037 NETTRAN_DUMMY_1038 MUX2_X1 
XU334 n1634 n1625 n484 n333 NETTRAN_DUMMY_1039 NETTRAN_DUMMY_1040 MUX2_X1 
XU333 n331 n327 addr[4] n332 NETTRAN_DUMMY_1041 NETTRAN_DUMMY_1042 MUX2_X1 
XU332 n330 n329 addr[2] n331 NETTRAN_DUMMY_1043 NETTRAN_DUMMY_1044 MUX2_X1 
XU331 n1625 n1612 n484 n330 NETTRAN_DUMMY_1045 NETTRAN_DUMMY_1046 MUX2_X1 
XU330 n328 n7 n484 n329 NETTRAN_DUMMY_1047 NETTRAN_DUMMY_1048 MUX2_X1 
XU328 n326 n325 addr[2] n327 NETTRAN_DUMMY_1049 NETTRAN_DUMMY_1050 MUX2_X1 
XU327 n1639 n8 addr[3] n326 NETTRAN_DUMMY_1051 NETTRAN_DUMMY_1052 MUX2_X1 
XU326 n1653 n451 n484 n325 NETTRAN_DUMMY_1053 NETTRAN_DUMMY_1054 MUX2_X1 
XU325 n323 n313 addr[7] n324 NETTRAN_DUMMY_1055 NETTRAN_DUMMY_1056 MUX2_X1 
XU324 n322 n318 addr[4] n323 NETTRAN_DUMMY_1057 NETTRAN_DUMMY_1058 MUX2_X1 
XU323 n321 n319 addr[2] n322 NETTRAN_DUMMY_1059 NETTRAN_DUMMY_1060 MUX2_X1 
XU322 n512 n320 n484 n321 NETTRAN_DUMMY_1061 NETTRAN_DUMMY_1062 MUX2_X1 
XU321 n5 addr[0] addr[5] n320 NETTRAN_DUMMY_1063 NETTRAN_DUMMY_1064 MUX2_X1 
XU320 n25 n51 n484 n319 NETTRAN_DUMMY_1065 NETTRAN_DUMMY_1066 MUX2_X1 
XU319 n315 n316 addr[2] n318 NETTRAN_DUMMY_1067 NETTRAN_DUMMY_1068 MUX2_X1 
XU317 n314 n1595 n484 n315 NETTRAN_DUMMY_1069 NETTRAN_DUMMY_1070 MUX2_X1 
XU316 n512 n1 addr[5] n314 NETTRAN_DUMMY_1071 NETTRAN_DUMMY_1072 MUX2_X1 
XU315 n312 n307 addr[4] n313 NETTRAN_DUMMY_1073 NETTRAN_DUMMY_1074 MUX2_X1 
XU314 n309 n310 addr[2] n312 NETTRAN_DUMMY_1075 NETTRAN_DUMMY_1076 MUX2_X1 
XU312 n1626 n308 n484 n309 NETTRAN_DUMMY_1077 NETTRAN_DUMMY_1078 MUX2_X1 
XU311 n1537 n9 addr[5] n308 NETTRAN_DUMMY_1079 NETTRAN_DUMMY_1080 MUX2_X1 
XU310 n306 n305 addr[2] n307 NETTRAN_DUMMY_1081 NETTRAN_DUMMY_1082 MUX2_X1 
XU308 n1599 n451 n484 n305 NETTRAN_DUMMY_1083 NETTRAN_DUMMY_1084 MUX2_X1 
XU307 n304 n289 addr[6] d[6] NETTRAN_DUMMY_1085 NETTRAN_DUMMY_1086 MUX2_X1 
XU306 n303 n296 addr[7] n304 NETTRAN_DUMMY_1087 NETTRAN_DUMMY_1088 MUX2_X1 
XU305 n302 n299 n460 n303 NETTRAN_DUMMY_1089 NETTRAN_DUMMY_1090 MUX2_X1 
XU304 n301 n300 IN0 n302 NETTRAN_DUMMY_1091 NETTRAN_DUMMY_1092 MUX2_X1 
XU303 n1612 n1661 n487 n301 NETTRAN_DUMMY_1093 NETTRAN_DUMMY_1094 MUX2_X1 
XU302 n1660 n1641 n487 n300 NETTRAN_DUMMY_1095 NETTRAN_DUMMY_1096 MUX2_X1 
XU301 n298 n297 IN0 n299 NETTRAN_DUMMY_1097 NETTRAN_DUMMY_1098 MUX2_X1 
XU299 n1610 n54 n487 n297 NETTRAN_DUMMY_1099 NETTRAN_DUMMY_1100 MUX2_X1 
XU298 n295 n292 n460 n296 NETTRAN_DUMMY_1101 NETTRAN_DUMMY_1102 MUX2_X1 
XU297 n294 n293 addr[2] n295 NETTRAN_DUMMY_1103 NETTRAN_DUMMY_1104 MUX2_X1 
XU296 n50 n35 addr[3] n294 NETTRAN_DUMMY_1105 NETTRAN_DUMMY_1106 MUX2_X1 
XU295 n1637 n16 addr[3] n293 NETTRAN_DUMMY_1107 NETTRAN_DUMMY_1108 MUX2_X1 
XU294 n291 n290 addr[2] n292 NETTRAN_DUMMY_1109 NETTRAN_DUMMY_1110 MUX2_X1 
XU293 n15 n1640 addr[3] n291 NETTRAN_DUMMY_1111 NETTRAN_DUMMY_1112 MUX2_X1 
XU292 n1660 n53 n487 n290 NETTRAN_DUMMY_1113 NETTRAN_DUMMY_1114 MUX2_X1 
XU291 n288 n281 addr[7] n289 NETTRAN_DUMMY_1115 NETTRAN_DUMMY_1116 MUX2_X1 
XU290 n287 n284 n460 n288 NETTRAN_DUMMY_1117 NETTRAN_DUMMY_1118 MUX2_X1 
XU289 n286 n285 IN0 n287 NETTRAN_DUMMY_1119 NETTRAN_DUMMY_1120 MUX2_X1 
XU288 n1633 n1641 n487 n286 NETTRAN_DUMMY_1121 NETTRAN_DUMMY_1122 MUX2_X1 
XU287 n21 n4 n487 n285 NETTRAN_DUMMY_1123 NETTRAN_DUMMY_1124 MUX2_X1 
XU286 n283 n282 IN0 n284 NETTRAN_DUMMY_1125 NETTRAN_DUMMY_1126 MUX2_X1 
XU285 n1659 n40 n487 n283 NETTRAN_DUMMY_1127 NETTRAN_DUMMY_1128 MUX2_X1 
XU284 n1594 n1622 n487 n282 NETTRAN_DUMMY_1129 NETTRAN_DUMMY_1130 MUX2_X1 
XU283 n280 n277 addr[4] n281 NETTRAN_DUMMY_1131 NETTRAN_DUMMY_1132 MUX2_X1 
XU282 n279 n278 addr[2] n280 NETTRAN_DUMMY_1133 NETTRAN_DUMMY_1134 MUX2_X1 
XU281 n1625 n1629 addr[3] n279 NETTRAN_DUMMY_1135 NETTRAN_DUMMY_1136 MUX2_X1 
XU280 n1647 n1594 addr[3] n278 NETTRAN_DUMMY_1137 NETTRAN_DUMMY_1138 MUX2_X1 
XU279 n1600 n276 n429 n277 NETTRAN_DUMMY_1139 NETTRAN_DUMMY_1140 MUX2_X1 
XU278 n1591 n1536 n492 n276 NETTRAN_DUMMY_1141 NETTRAN_DUMMY_1142 MUX2_X1 
XU277 n275 n257 addr[6] d[5] NETTRAN_DUMMY_1143 NETTRAN_DUMMY_1144 MUX2_X1 
XU276 n274 n265 n460 n275 NETTRAN_DUMMY_1145 NETTRAN_DUMMY_1146 MUX2_X1 
XU275 n273 n268 addr[2] n274 NETTRAN_DUMMY_1147 NETTRAN_DUMMY_1148 MUX2_X1 
XU274 n272 n270 n487 n273 NETTRAN_DUMMY_1149 NETTRAN_DUMMY_1150 MUX2_X1 
XU619 n533 n1520 n515 n608 NETTRAN_DUMMY_1151 NETTRAN_DUMMY_1152 MUX2_X1 
XU617 n1522 n492 n509 n606 NETTRAN_DUMMY_1153 NETTRAN_DUMMY_1154 MUX2_X1 
XU616 n1526 n1522 n515 n605 NETTRAN_DUMMY_1155 NETTRAN_DUMMY_1156 MUX2_X1 
XU614 n517 n1522 n509 n603 NETTRAN_DUMMY_1157 NETTRAN_DUMMY_1158 MUX2_X1 
XU613 n488 n492 n515 n602 NETTRAN_DUMMY_1159 NETTRAN_DUMMY_1160 MUX2_X1 
XU612 n1526 n488 n515 n601 NETTRAN_DUMMY_1161 NETTRAN_DUMMY_1162 MUX2_X1 
XU610 n488 n528 n509 n599 NETTRAN_DUMMY_1163 NETTRAN_DUMMY_1164 MUX2_X1 
XU609 n492 n480 n513 n598 NETTRAN_DUMMY_1165 NETTRAN_DUMMY_1166 MUX2_X1 
XU607 n1318 n492 n515 n596 NETTRAN_DUMMY_1167 NETTRAN_DUMMY_1168 MUX2_X1 
XU606 n526 n492 n509 n595 NETTRAN_DUMMY_1169 NETTRAN_DUMMY_1170 MUX2_X1 
XU605 n493 n517 n509 n594 NETTRAN_DUMMY_1171 NETTRAN_DUMMY_1172 MUX2_X1 
XU602 n1318 n1522 n515 n591 NETTRAN_DUMMY_1173 NETTRAN_DUMMY_1174 MUX2_X1 
XU601 n517 n515 n590 NETTRAN_DUMMY_1175 NETTRAN_DUMMY_1176 XOR2_X1 
XU600 n492 n1526 n509 n589 NETTRAN_DUMMY_1177 NETTRAN_DUMMY_1178 MUX2_X1 
XU599 IN1 n526 n515 n588 NETTRAN_DUMMY_1179 NETTRAN_DUMMY_1180 MUX2_X1 
XU597 n517 n488 n509 n586 NETTRAN_DUMMY_1181 NETTRAN_DUMMY_1182 MUX2_X1 
XU596 n1525 n1526 n515 n585 NETTRAN_DUMMY_1183 NETTRAN_DUMMY_1184 MUX2_X1 
XU595 n1525 n492 n509 n584 NETTRAN_DUMMY_1185 NETTRAN_DUMMY_1186 MUX2_X1 
XU594 n533 n492 n515 n583 NETTRAN_DUMMY_1187 NETTRAN_DUMMY_1188 MUX2_X1 
XU590 n488 n513 n579 NETTRAN_DUMMY_1189 NETTRAN_DUMMY_1190 XOR2_X1 
XU589 n520 IN1 n515 n578 NETTRAN_DUMMY_1191 NETTRAN_DUMMY_1192 MUX2_X1 
XU588 n520 n526 n509 n577 NETTRAN_DUMMY_1193 NETTRAN_DUMMY_1194 MUX2_X1 
XU587 n492 n1520 n515 n576 NETTRAN_DUMMY_1195 NETTRAN_DUMMY_1196 MUX2_X1 
XU586 n517 n492 n515 n575 NETTRAN_DUMMY_1197 NETTRAN_DUMMY_1198 MUX2_X1 
XU584 n488 n533 n515 n573 NETTRAN_DUMMY_1199 NETTRAN_DUMMY_1200 MUX2_X1 
XU583 n480 n520 n513 n547 NETTRAN_DUMMY_1201 NETTRAN_DUMMY_1202 MUX2_X1 
XU582 n1520 n1526 n515 n572 NETTRAN_DUMMY_1203 NETTRAN_DUMMY_1204 MUX2_X1 
XU581 n1522 IN1 n515 n571 NETTRAN_DUMMY_1205 NETTRAN_DUMMY_1206 MUX2_X1 
XU580 n492 n528 n515 n570 NETTRAN_DUMMY_1207 NETTRAN_DUMMY_1208 MUX2_X1 
XU578 n449 n468 n568 NETTRAN_DUMMY_1209 NETTRAN_DUMMY_1210 XOR2_X1 
XU577 n488 n526 n515 n567 NETTRAN_DUMMY_1211 NETTRAN_DUMMY_1212 MUX2_X1 
XU576 n1526 n1318 n515 n566 NETTRAN_DUMMY_1213 NETTRAN_DUMMY_1214 MUX2_X1 
XU575 n533 n526 n509 n565 NETTRAN_DUMMY_1215 NETTRAN_DUMMY_1216 MUX2_X1 
XU574 n492 n1522 n515 n564 NETTRAN_DUMMY_1217 NETTRAN_DUMMY_1218 MUX2_X1 
XU573 n1522 n517 n509 n563 NETTRAN_DUMMY_1219 NETTRAN_DUMMY_1220 MUX2_X1 
XU572 IN1 n492 n515 n562 NETTRAN_DUMMY_1221 NETTRAN_DUMMY_1222 MUX2_X1 
XU571 n512 n1522 n561 NETTRAN_DUMMY_1223 NETTRAN_DUMMY_1224 XOR2_X1 
XU569 n528 n517 n509 n559 NETTRAN_DUMMY_1225 NETTRAN_DUMMY_1226 MUX2_X1 
XU567 n533 IN1 n515 n557 NETTRAN_DUMMY_1227 NETTRAN_DUMMY_1228 MUX2_X1 
XU566 n528 n520 n509 n556 NETTRAN_DUMMY_1229 NETTRAN_DUMMY_1230 MUX2_X1 
XU564 n488 n1522 n509 n554 NETTRAN_DUMMY_1231 NETTRAN_DUMMY_1232 MUX2_X1 
XU563 n1318 n1525 n515 n553 NETTRAN_DUMMY_1233 NETTRAN_DUMMY_1234 MUX2_X1 
XU557 n1520 n533 n509 n550 NETTRAN_DUMMY_1235 NETTRAN_DUMMY_1236 MUX2_X1 
XU556 n493 n1318 n509 n549 NETTRAN_DUMMY_1237 NETTRAN_DUMMY_1238 MUX2_X1 
XU554 n488 n492 n533 NETTRAN_DUMMY_1239 NETTRAN_DUMMY_1240 XOR2_X1 
XU439 n1614 n1610 n487 n402 NETTRAN_DUMMY_1241 NETTRAN_DUMMY_1242 MUX2_X1 
XU438 n426 n461 n487 n403 NETTRAN_DUMMY_1243 NETTRAN_DUMMY_1244 MUX2_X1 
XU436 addr[0] n9 n448 n425 NETTRAN_DUMMY_1245 NETTRAN_DUMMY_1246 MUX2_X1 
XU435 n406 n13 n480 n347 NETTRAN_DUMMY_1247 NETTRAN_DUMMY_1248 MUX2_X1 
XU434 addr[0] n1 n448 n424 NETTRAN_DUMMY_1249 NETTRAN_DUMMY_1250 MUX2_X1 
XU433 n501 n1 n448 n423 NETTRAN_DUMMY_1251 NETTRAN_DUMMY_1252 MUX2_X1 
XU432 n1540 n1531 addr[5] n422 NETTRAN_DUMMY_1253 NETTRAN_DUMMY_1254 MUX2_X1 
XU431 n5 n2 addr[5] n421 NETTRAN_DUMMY_1255 NETTRAN_DUMMY_1256 MUX2_X1 
XU430 addr[1] n2 addr[5] n420 NETTRAN_DUMMY_1257 NETTRAN_DUMMY_1258 MUX2_X1 
XU429 n41 n43 addr[2] n223 NETTRAN_DUMMY_1259 NETTRAN_DUMMY_1260 MUX2_X1 
XU428 n1646 n449 n480 n201 NETTRAN_DUMMY_1261 NETTRAN_DUMMY_1262 MUX2_X1 
XU427 n1540 addr[1] addr[5] n419 NETTRAN_DUMMY_1263 NETTRAN_DUMMY_1264 MUX2_X1 
XU426 n501 n1540 n448 n418 NETTRAN_DUMMY_1265 NETTRAN_DUMMY_1266 MUX2_X1 
XU425 n455 n38 IN0 n417 NETTRAN_DUMMY_1267 NETTRAN_DUMMY_1268 MUX2_X1 
XU424 n501 n6 n448 n416 NETTRAN_DUMMY_1269 NETTRAN_DUMMY_1270 MUX2_X1 
XU423 n1537 addr[1] addr[5] n415 NETTRAN_DUMMY_1271 NETTRAN_DUMMY_1272 MUX2_X1 
XU422 n2 n1531 n448 n414 NETTRAN_DUMMY_1273 NETTRAN_DUMMY_1274 MUX2_X1 
XU421 n512 n9 n448 n413 NETTRAN_DUMMY_1275 NETTRAN_DUMMY_1276 MUX2_X1 
XU420 n1623 n407 n460 n412 NETTRAN_DUMMY_1277 NETTRAN_DUMMY_1278 MUX2_X1 
XU407 n9 n1527 addr[5] n221 NETTRAN_DUMMY_1279 NETTRAN_DUMMY_1280 MUX2_X1 
XU406 n405 n389 addr[6] d[9] NETTRAN_DUMMY_1281 NETTRAN_DUMMY_1282 MUX2_X1 
XU405 n404 n397 addr[7] n405 NETTRAN_DUMMY_1283 NETTRAN_DUMMY_1284 MUX2_X1 
XU404 n400 n401 IN0 n404 NETTRAN_DUMMY_1285 NETTRAN_DUMMY_1286 MUX2_X1 
XU402 n399 n398 n487 n400 NETTRAN_DUMMY_1287 NETTRAN_DUMMY_1288 MUX2_X1 
XU401 n1 n1644 n460 n399 NETTRAN_DUMMY_1289 NETTRAN_DUMMY_1290 MUX2_X1 
XU400 n41 n1662 n460 n398 NETTRAN_DUMMY_1291 NETTRAN_DUMMY_1292 MUX2_X1 
XU399 n396 n392 IN0 n397 NETTRAN_DUMMY_1293 NETTRAN_DUMMY_1294 MUX2_X1 
XU398 n395 n393 n484 n396 NETTRAN_DUMMY_1295 NETTRAN_DUMMY_1296 MUX2_X1 
XU397 n1654 n394 addr[4] n395 NETTRAN_DUMMY_1297 NETTRAN_DUMMY_1298 MUX2_X1 
XU396 n512 n1524 addr[5] n394 NETTRAN_DUMMY_1299 NETTRAN_DUMMY_1300 MUX2_X1 
XU395 n52 n1657 addr[4] n393 NETTRAN_DUMMY_1301 NETTRAN_DUMMY_1302 MUX2_X1 
XU394 n391 n390 n487 n392 NETTRAN_DUMMY_1303 NETTRAN_DUMMY_1304 MUX2_X1 
XU393 n55 n59 n460 n391 NETTRAN_DUMMY_1305 NETTRAN_DUMMY_1306 MUX2_X1 
XU392 n1662 n1638 n460 n390 NETTRAN_DUMMY_1307 NETTRAN_DUMMY_1308 MUX2_X1 
XU391 n388 n381 addr[7] n389 NETTRAN_DUMMY_1309 NETTRAN_DUMMY_1310 MUX2_X1 
XU390 n387 n384 addr[2] n388 NETTRAN_DUMMY_1311 NETTRAN_DUMMY_1312 MUX2_X1 
XU389 n386 n385 n487 n387 NETTRAN_DUMMY_1313 NETTRAN_DUMMY_1314 MUX2_X1 
XU388 n57 n1642 n460 n386 NETTRAN_DUMMY_1315 NETTRAN_DUMMY_1316 MUX2_X1 
XU387 n1536 n1649 n460 n385 NETTRAN_DUMMY_1317 NETTRAN_DUMMY_1318 MUX2_X1 
XU386 n383 n382 n487 n384 NETTRAN_DUMMY_1319 NETTRAN_DUMMY_1320 MUX2_X1 
XU385 n1616 n1659 n460 n383 NETTRAN_DUMMY_1321 NETTRAN_DUMMY_1322 MUX2_X1 
XU384 n49 n1631 n460 n382 NETTRAN_DUMMY_1323 NETTRAN_DUMMY_1324 MUX2_X1 
XU383 n380 n377 addr[2] n381 NETTRAN_DUMMY_1325 NETTRAN_DUMMY_1326 MUX2_X1 
XU382 n379 n378 n487 n380 NETTRAN_DUMMY_1327 NETTRAN_DUMMY_1328 MUX2_X1 
XU380 n1595 n1536 n460 n378 NETTRAN_DUMMY_1329 NETTRAN_DUMMY_1330 MUX2_X1 
XU379 n1604 n376 n487 n377 NETTRAN_DUMMY_1331 NETTRAN_DUMMY_1332 MUX2_X1 
XU378 n1597 n1593 n460 n376 NETTRAN_DUMMY_1333 NETTRAN_DUMMY_1334 MUX2_X1 
XU377 n375 n357 addr[6] d[8] NETTRAN_DUMMY_1335 NETTRAN_DUMMY_1336 MUX2_X1 
XU723 n1501 n537 n445 n709 NETTRAN_DUMMY_1337 NETTRAN_DUMMY_1338 MUX2_X1 
XU722 n708 n696 n433 d[11] NETTRAN_DUMMY_1339 NETTRAN_DUMMY_1340 MUX2_X1 
XU721 n707 n700 n439 n708 NETTRAN_DUMMY_1341 NETTRAN_DUMMY_1342 MUX2_X1 
XU720 n706 n703 n503 n707 NETTRAN_DUMMY_1343 NETTRAN_DUMMY_1344 MUX2_X1 
XU719 n705 n704 n452 n706 NETTRAN_DUMMY_1345 NETTRAN_DUMMY_1346 MUX2_X1 
XU718 n604 n538 n473 n705 NETTRAN_DUMMY_1347 NETTRAN_DUMMY_1348 MUX2_X1 
XU717 n1846 n1776 n462 n704 NETTRAN_DUMMY_1349 NETTRAN_DUMMY_1350 MUX2_X1 
XU716 n702 n701 n452 n703 NETTRAN_DUMMY_1351 NETTRAN_DUMMY_1352 MUX2_X1 
XU715 n1528 n493 n473 n702 NETTRAN_DUMMY_1353 NETTRAN_DUMMY_1354 MUX2_X1 
XU714 n1796 n1833 n473 n701 NETTRAN_DUMMY_1355 NETTRAN_DUMMY_1356 MUX2_X1 
XU713 n699 n697 n503 n700 NETTRAN_DUMMY_1357 NETTRAN_DUMMY_1358 MUX2_X1 
XU712 n698 n631 n452 n699 NETTRAN_DUMMY_1359 NETTRAN_DUMMY_1360 MUX2_X1 
XU711 n1787 n1318 n462 n698 NETTRAN_DUMMY_1361 NETTRAN_DUMMY_1362 MUX2_X1 
XU710 n630 n574 n452 n697 NETTRAN_DUMMY_1363 NETTRAN_DUMMY_1364 MUX2_X1 
XU709 n695 n691 n439 n696 NETTRAN_DUMMY_1365 NETTRAN_DUMMY_1366 MUX2_X1 
XU708 n693 n694 n503 n695 NETTRAN_DUMMY_1367 NETTRAN_DUMMY_1368 MUX2_X1 
XU706 n1670 n692 n452 n693 NETTRAN_DUMMY_1369 NETTRAN_DUMMY_1370 MUX2_X1 
XU704 n690 n1663 n503 n691 NETTRAN_DUMMY_1371 NETTRAN_DUMMY_1372 MUX2_X1 
XU703 n689 n1665 n452 n690 NETTRAN_DUMMY_1373 NETTRAN_DUMMY_1374 MUX2_X1 
XU701 n688 n673 n433 d[10] NETTRAN_DUMMY_1375 NETTRAN_DUMMY_1376 MUX2_X1 
XU700 n687 n680 n442 n688 NETTRAN_DUMMY_1377 NETTRAN_DUMMY_1378 MUX2_X1 
XU699 n686 n683 n503 n687 NETTRAN_DUMMY_1379 NETTRAN_DUMMY_1380 MUX2_X1 
XU698 n685 n684 n452 n686 NETTRAN_DUMMY_1381 NETTRAN_DUMMY_1382 MUX2_X1 
XU697 n517 n1774 n473 n685 NETTRAN_DUMMY_1383 NETTRAN_DUMMY_1384 MUX2_X1 
XU696 n522 n1848 n473 n684 NETTRAN_DUMMY_1385 NETTRAN_DUMMY_1386 MUX2_X1 
XU695 n682 n681 n452 n683 NETTRAN_DUMMY_1387 NETTRAN_DUMMY_1388 MUX2_X1 
XU694 n1811 n1333 n473 n682 NETTRAN_DUMMY_1389 NETTRAN_DUMMY_1390 MUX2_X1 
XU693 n1533 n1775 n475 n681 NETTRAN_DUMMY_1391 NETTRAN_DUMMY_1392 MUX2_X1 
XU692 n679 n676 n503 n680 NETTRAN_DUMMY_1393 NETTRAN_DUMMY_1394 MUX2_X1 
XU691 n678 n677 n452 n679 NETTRAN_DUMMY_1395 NETTRAN_DUMMY_1396 MUX2_X1 
XU690 n629 n533 n473 n678 NETTRAN_DUMMY_1397 NETTRAN_DUMMY_1398 MUX2_X1 
XU689 n1534 n1789 n473 n677 NETTRAN_DUMMY_1399 NETTRAN_DUMMY_1400 MUX2_X1 
XU688 n675 n674 n452 n676 NETTRAN_DUMMY_1401 NETTRAN_DUMMY_1402 MUX2_X1 
XU686 n1318 n535 n473 n674 NETTRAN_DUMMY_1403 NETTRAN_DUMMY_1404 MUX2_X1 
XU685 n672 n666 n445 n673 NETTRAN_DUMMY_1405 NETTRAN_DUMMY_1406 MUX2_X1 
XU684 n671 n668 n503 n672 NETTRAN_DUMMY_1407 NETTRAN_DUMMY_1408 MUX2_X1 
XU683 n670 n669 n452 n671 NETTRAN_DUMMY_1409 NETTRAN_DUMMY_1410 MUX2_X1 
XU682 n532 n1535 n473 n670 NETTRAN_DUMMY_1411 NETTRAN_DUMMY_1412 MUX2_X1 
XU681 n1541 n524 n473 n669 NETTRAN_DUMMY_1413 NETTRAN_DUMMY_1414 MUX2_X1 
XU680 n534 n667 n452 n668 NETTRAN_DUMMY_1415 NETTRAN_DUMMY_1416 MUX2_X1 
XU679 n536 n513 n473 n667 NETTRAN_DUMMY_1417 NETTRAN_DUMMY_1418 MUX2_X1 
XU678 n665 n1663 n497 n666 NETTRAN_DUMMY_1419 NETTRAN_DUMMY_1420 MUX2_X1 
XU676 n1545 n1318 n448 n664 NETTRAN_DUMMY_1421 NETTRAN_DUMMY_1422 MUX2_X1 
XU675 n663 n648 n433 d[0] NETTRAN_DUMMY_1423 NETTRAN_DUMMY_1424 MUX2_X1 
XU674 n662 n655 n452 n663 NETTRAN_DUMMY_1425 NETTRAN_DUMMY_1426 MUX2_X1 
XU673 n661 n658 n497 n662 NETTRAN_DUMMY_1427 NETTRAN_DUMMY_1428 MUX2_X1 
XU672 n659 n660 n458 n661 NETTRAN_DUMMY_1429 NETTRAN_DUMMY_1430 MUX2_X1 
XU670 n518 n1544 n443 n659 NETTRAN_DUMMY_1431 NETTRAN_DUMMY_1432 MUX2_X1 
XU669 n657 n656 n473 n658 NETTRAN_DUMMY_1433 NETTRAN_DUMMY_1434 MUX2_X1 
XU668 n1822 n1790 n443 n657 NETTRAN_DUMMY_1435 NETTRAN_DUMMY_1436 MUX2_X1 
XU667 n1526 n1501 n442 n656 NETTRAN_DUMMY_1437 NETTRAN_DUMMY_1438 MUX2_X1 
XU666 n654 n651 n497 n655 NETTRAN_DUMMY_1439 NETTRAN_DUMMY_1440 MUX2_X1 
XU665 n653 n652 n473 n654 NETTRAN_DUMMY_1441 NETTRAN_DUMMY_1442 MUX2_X1 
XU664 n628 n524 n442 n653 NETTRAN_DUMMY_1443 NETTRAN_DUMMY_1444 MUX2_X1 
XU663 n527 n529 n445 n652 NETTRAN_DUMMY_1445 NETTRAN_DUMMY_1446 MUX2_X1 
XU662 n650 n649 n473 n651 NETTRAN_DUMMY_1447 NETTRAN_DUMMY_1448 MUX2_X1 
XU661 n526 n1499 n442 n650 NETTRAN_DUMMY_1449 NETTRAN_DUMMY_1450 MUX2_X1 
XU660 n1501 n1754 n442 n649 NETTRAN_DUMMY_1451 NETTRAN_DUMMY_1452 MUX2_X1 
XU659 n647 n640 n452 n648 NETTRAN_DUMMY_1453 NETTRAN_DUMMY_1454 MUX2_X1 
XU658 n646 n643 n507 n647 NETTRAN_DUMMY_1455 NETTRAN_DUMMY_1456 MUX2_X1 
XU657 n645 n644 n475 n646 NETTRAN_DUMMY_1457 NETTRAN_DUMMY_1458 MUX2_X1 
XU656 n1674 n1772 n443 n645 NETTRAN_DUMMY_1459 NETTRAN_DUMMY_1460 MUX2_X1 
XU655 n1855 n509 n443 n644 NETTRAN_DUMMY_1461 NETTRAN_DUMMY_1462 MUX2_X1 
XU654 n642 n641 n475 n643 NETTRAN_DUMMY_1463 NETTRAN_DUMMY_1464 MUX2_X1 
XU653 n521 n1835 n443 n642 NETTRAN_DUMMY_1465 NETTRAN_DUMMY_1466 MUX2_X1 
XU652 n550 n530 n443 n641 NETTRAN_DUMMY_1467 NETTRAN_DUMMY_1468 MUX2_X1 
XU651 n639 n636 n503 n640 NETTRAN_DUMMY_1469 NETTRAN_DUMMY_1470 MUX2_X1 
XU650 n637 n638 n473 n639 NETTRAN_DUMMY_1471 NETTRAN_DUMMY_1472 MUX2_X1 
XU648 n1773 n1789 n439 n637 NETTRAN_DUMMY_1473 NETTRAN_DUMMY_1474 MUX2_X1 
XU647 n634 n635 n473 n636 NETTRAN_DUMMY_1475 NETTRAN_DUMMY_1476 MUX2_X1 
XU645 n1808 n1765 n442 n634 NETTRAN_DUMMY_1477 NETTRAN_DUMMY_1478 MUX2_X1 
XU644 n517 n464 n633 NETTRAN_DUMMY_1479 NETTRAN_DUMMY_1480 XOR2_X1 
XU643 n461 n513 n632 NETTRAN_DUMMY_1481 NETTRAN_DUMMY_1482 XOR2_X1 
XU642 n461 n1538 n631 NETTRAN_DUMMY_1483 NETTRAN_DUMMY_1484 XOR2_X1 
XU641 n539 n473 n630 NETTRAN_DUMMY_1485 NETTRAN_DUMMY_1486 XOR2_X1 
XU640 n493 n509 n629 NETTRAN_DUMMY_1487 NETTRAN_DUMMY_1488 XOR2_X1 
XU639 n520 n513 n628 NETTRAN_DUMMY_1489 NETTRAN_DUMMY_1490 XOR2_X1 
XU638 n526 n513 n627 NETTRAN_DUMMY_1491 NETTRAN_DUMMY_1492 XOR2_X1 
XU637 n528 n515 n626 NETTRAN_DUMMY_1493 NETTRAN_DUMMY_1494 XOR2_X1 
XU634 n512 n1501 n473 n623 NETTRAN_DUMMY_1495 NETTRAN_DUMMY_1496 MUX2_X1 
XU633 n1318 n480 n509 n622 NETTRAN_DUMMY_1497 NETTRAN_DUMMY_1498 MUX2_X1 
XU632 n1525 n488 n509 n621 NETTRAN_DUMMY_1499 NETTRAN_DUMMY_1500 MUX2_X1 
XU631 n1520 n492 n509 n620 NETTRAN_DUMMY_1501 NETTRAN_DUMMY_1502 MUX2_X1 
XU630 n480 n1318 n513 n619 NETTRAN_DUMMY_1503 NETTRAN_DUMMY_1504 MUX2_X1 
XU629 n488 n1525 n515 n618 NETTRAN_DUMMY_1505 NETTRAN_DUMMY_1506 MUX2_X1 
XU628 n493 n1525 n515 n617 NETTRAN_DUMMY_1507 NETTRAN_DUMMY_1508 MUX2_X1 
XU626 n493 n1522 n509 n615 NETTRAN_DUMMY_1509 NETTRAN_DUMMY_1510 MUX2_X1 
XU625 n1318 n493 n509 n614 NETTRAN_DUMMY_1511 NETTRAN_DUMMY_1512 MUX2_X1 
XU624 n528 n492 n515 n613 NETTRAN_DUMMY_1513 NETTRAN_DUMMY_1514 MUX2_X1 
XU623 n526 n488 n509 n612 NETTRAN_DUMMY_1515 NETTRAN_DUMMY_1516 MUX2_X1 
XU622 n520 n528 n509 n611 NETTRAN_DUMMY_1517 NETTRAN_DUMMY_1518 MUX2_X1 
XU621 n533 n520 n509 n610 NETTRAN_DUMMY_1519 NETTRAN_DUMMY_1520 MUX2_X1 
XU620 n1525 n1520 n509 n609 NETTRAN_DUMMY_1521 NETTRAN_DUMMY_1522 MUX2_X1 
XU835 n820 n805 n433 d[18] NETTRAN_DUMMY_1523 NETTRAN_DUMMY_1524 MUX2_X1 
XU834 n819 n812 n455 n820 NETTRAN_DUMMY_1525 NETTRAN_DUMMY_1526 MUX2_X1 
XU833 n818 n815 n495 n819 NETTRAN_DUMMY_1527 NETTRAN_DUMMY_1528 MUX2_X1 
XU832 n1756 n816 n458 n818 NETTRAN_DUMMY_1529 NETTRAN_DUMMY_1530 MUX2_X1 
XU830 n814 n813 n471 n815 NETTRAN_DUMMY_1531 NETTRAN_DUMMY_1532 MUX2_X1 
XU829 n1838 n1760 n443 n814 NETTRAN_DUMMY_1533 NETTRAN_DUMMY_1534 MUX2_X1 
XU828 n589 n1543 n443 n813 NETTRAN_DUMMY_1535 NETTRAN_DUMMY_1536 MUX2_X1 
XU827 n811 n808 n495 n812 NETTRAN_DUMMY_1537 NETTRAN_DUMMY_1538 MUX2_X1 
XU826 n810 n809 n471 n811 NETTRAN_DUMMY_1539 NETTRAN_DUMMY_1540 MUX2_X1 
XU825 n1743 n1842 n443 n810 NETTRAN_DUMMY_1541 NETTRAN_DUMMY_1542 MUX2_X1 
XU824 n531 n1534 n443 n809 NETTRAN_DUMMY_1543 NETTRAN_DUMMY_1544 MUX2_X1 
XU823 n806 n807 n471 n808 NETTRAN_DUMMY_1545 NETTRAN_DUMMY_1546 MUX2_X1 
XU821 n532 n572 n443 n806 NETTRAN_DUMMY_1547 NETTRAN_DUMMY_1548 MUX2_X1 
XU820 n804 n797 n455 n805 NETTRAN_DUMMY_1549 NETTRAN_DUMMY_1550 MUX2_X1 
XU819 n803 n800 n495 n804 NETTRAN_DUMMY_1551 NETTRAN_DUMMY_1552 MUX2_X1 
XU818 n802 n801 n471 n803 NETTRAN_DUMMY_1553 NETTRAN_DUMMY_1554 MUX2_X1 
XU817 n586 n1804 n443 n802 NETTRAN_DUMMY_1555 NETTRAN_DUMMY_1556 MUX2_X1 
XU816 n1824 n1774 n443 n801 NETTRAN_DUMMY_1557 NETTRAN_DUMMY_1558 MUX2_X1 
XU815 n799 n798 n471 n800 NETTRAN_DUMMY_1559 NETTRAN_DUMMY_1560 MUX2_X1 
XU814 n1797 n1760 n443 n799 NETTRAN_DUMMY_1561 NETTRAN_DUMMY_1562 MUX2_X1 
XU813 n1795 n1535 n443 n798 NETTRAN_DUMMY_1563 NETTRAN_DUMMY_1564 MUX2_X1 
XU812 n795 n796 n495 n797 NETTRAN_DUMMY_1565 NETTRAN_DUMMY_1566 MUX2_X1 
XU810 n793 n794 n471 n795 NETTRAN_DUMMY_1567 NETTRAN_DUMMY_1568 MUX2_X1 
XU808 n1811 n555 n443 n793 NETTRAN_DUMMY_1569 NETTRAN_DUMMY_1570 MUX2_X1 
XU807 n1500 n539 n458 n792 NETTRAN_DUMMY_1571 NETTRAN_DUMMY_1572 MUX2_X1 
XU806 n597 n445 n458 n791 NETTRAN_DUMMY_1573 NETTRAN_DUMMY_1574 MUX2_X1 
XU805 n790 n774 n433 d[17] NETTRAN_DUMMY_1575 NETTRAN_DUMMY_1576 MUX2_X1 
XU804 n789 n782 n445 n790 NETTRAN_DUMMY_1577 NETTRAN_DUMMY_1578 MUX2_X1 
XU803 n788 n785 n455 n789 NETTRAN_DUMMY_1579 NETTRAN_DUMMY_1580 MUX2_X1 
XU802 n787 n786 n495 n788 NETTRAN_DUMMY_1581 NETTRAN_DUMMY_1582 MUX2_X1 
XU801 n569 n1838 n471 n787 NETTRAN_DUMMY_1583 NETTRAN_DUMMY_1584 MUX2_X1 
XU800 n1523 n540 n471 n786 NETTRAN_DUMMY_1585 NETTRAN_DUMMY_1586 MUX2_X1 
XU799 n784 n783 n495 n785 NETTRAN_DUMMY_1587 NETTRAN_DUMMY_1588 MUX2_X1 
XU798 n1741 n541 n471 n784 NETTRAN_DUMMY_1589 NETTRAN_DUMMY_1590 MUX2_X1 
XU797 n1742 n1762 n471 n783 NETTRAN_DUMMY_1591 NETTRAN_DUMMY_1592 MUX2_X1 
XU796 n781 n778 n455 n782 NETTRAN_DUMMY_1593 NETTRAN_DUMMY_1594 MUX2_X1 
XU795 n780 n779 n495 n781 NETTRAN_DUMMY_1595 NETTRAN_DUMMY_1596 MUX2_X1 
XU794 n1743 n627 n458 n780 NETTRAN_DUMMY_1597 NETTRAN_DUMMY_1598 MUX2_X1 
XU793 n1756 n1839 n458 n779 NETTRAN_DUMMY_1599 NETTRAN_DUMMY_1600 MUX2_X1 
XU792 n777 n775 n495 n778 NETTRAN_DUMMY_1601 NETTRAN_DUMMY_1602 MUX2_X1 
XU791 n1539 n776 n458 n777 NETTRAN_DUMMY_1603 NETTRAN_DUMMY_1604 MUX2_X1 
XU789 n1756 n1805 n458 n775 NETTRAN_DUMMY_1605 NETTRAN_DUMMY_1606 MUX2_X1 
XU788 n773 n766 n445 n774 NETTRAN_DUMMY_1607 NETTRAN_DUMMY_1608 MUX2_X1 
XU787 n772 n769 n455 n773 NETTRAN_DUMMY_1609 NETTRAN_DUMMY_1610 MUX2_X1 
XU786 n771 n770 n495 n772 NETTRAN_DUMMY_1611 NETTRAN_DUMMY_1612 MUX2_X1 
XU785 n1797 n539 n458 n771 NETTRAN_DUMMY_1613 NETTRAN_DUMMY_1614 MUX2_X1 
XU784 n1756 n573 n458 n770 NETTRAN_DUMMY_1615 NETTRAN_DUMMY_1616 MUX2_X1 
XU783 n768 n767 n507 n769 NETTRAN_DUMMY_1617 NETTRAN_DUMMY_1618 MUX2_X1 
XU782 n1761 n1777 n475 n768 NETTRAN_DUMMY_1619 NETTRAN_DUMMY_1620 MUX2_X1 
XU781 n1744 n1791 n475 n767 NETTRAN_DUMMY_1621 NETTRAN_DUMMY_1622 MUX2_X1 
XU780 n763 n764 n455 n766 NETTRAN_DUMMY_1623 NETTRAN_DUMMY_1624 MUX2_X1 
XU778 n762 n761 n495 n763 NETTRAN_DUMMY_1625 NETTRAN_DUMMY_1626 MUX2_X1 
XU777 n512 n1352 n458 n762 NETTRAN_DUMMY_1627 NETTRAN_DUMMY_1628 MUX2_X1 
XU776 n760 n1838 n458 n761 NETTRAN_DUMMY_1629 NETTRAN_DUMMY_1630 MUX2_X1 
XU774 n757 n758 n433 d[14] NETTRAN_DUMMY_1631 NETTRAN_DUMMY_1632 MUX2_X1 
XU772 n756 n752 n503 n757 NETTRAN_DUMMY_1633 NETTRAN_DUMMY_1634 MUX2_X1 
XU771 n755 n753 n442 n756 NETTRAN_DUMMY_1635 NETTRAN_DUMMY_1636 MUX2_X1 
XU770 n754 n632 n452 n755 NETTRAN_DUMMY_1637 NETTRAN_DUMMY_1638 MUX2_X1 
XU769 n577 n1849 n473 n754 NETTRAN_DUMMY_1639 NETTRAN_DUMMY_1640 MUX2_X1 
XU768 n513 n1671 n452 n753 NETTRAN_DUMMY_1641 NETTRAN_DUMMY_1642 MUX2_X1 
XU767 n751 n1663 n445 n752 NETTRAN_DUMMY_1643 NETTRAN_DUMMY_1644 MUX2_X1 
XU766 n1670 n750 n452 n751 NETTRAN_DUMMY_1645 NETTRAN_DUMMY_1646 MUX2_X1 
XU764 n749 n737 n433 d[13] NETTRAN_DUMMY_1647 NETTRAN_DUMMY_1648 MUX2_X1 
XU763 n748 n741 n445 n749 NETTRAN_DUMMY_1649 NETTRAN_DUMMY_1650 MUX2_X1 
XU762 n747 n744 n448 n748 NETTRAN_DUMMY_1651 NETTRAN_DUMMY_1652 MUX2_X1 
XU761 n746 n745 n468 n747 NETTRAN_DUMMY_1653 NETTRAN_DUMMY_1654 MUX2_X1 
XU760 n1832 n577 n497 n746 NETTRAN_DUMMY_1655 NETTRAN_DUMMY_1656 MUX2_X1 
XU759 n547 n1812 n497 n745 NETTRAN_DUMMY_1657 NETTRAN_DUMMY_1658 MUX2_X1 
XU758 n743 n742 n468 n744 NETTRAN_DUMMY_1659 NETTRAN_DUMMY_1660 MUX2_X1 
XU755 n739 n740 n452 n741 NETTRAN_DUMMY_1661 NETTRAN_DUMMY_1662 MUX2_X1 
XU753 n738 n513 n497 n739 NETTRAN_DUMMY_1663 NETTRAN_DUMMY_1664 MUX2_X1 
XU752 n581 n1528 n473 n738 NETTRAN_DUMMY_1665 NETTRAN_DUMMY_1666 MUX2_X1 
XU751 n736 n735 n439 n737 NETTRAN_DUMMY_1667 NETTRAN_DUMMY_1668 MUX2_X1 
XU749 n733 n732 n448 n735 NETTRAN_DUMMY_1669 NETTRAN_DUMMY_1670 MUX2_X1 
XU746 n531 n1318 n497 n731 NETTRAN_DUMMY_1671 NETTRAN_DUMMY_1672 MUX2_X1 
XU745 n730 n715 n433 d[12] NETTRAN_DUMMY_1673 NETTRAN_DUMMY_1674 MUX2_X1 
XU744 n729 n722 n497 n730 NETTRAN_DUMMY_1675 NETTRAN_DUMMY_1676 MUX2_X1 
XU743 n728 n725 n455 n729 NETTRAN_DUMMY_1677 NETTRAN_DUMMY_1678 MUX2_X1 
XU742 n727 n726 n458 n728 NETTRAN_DUMMY_1679 NETTRAN_DUMMY_1680 MUX2_X1 
XU741 n1763 n1535 n443 n727 NETTRAN_DUMMY_1681 NETTRAN_DUMMY_1682 MUX2_X1 
XU740 n1839 n628 n445 n726 NETTRAN_DUMMY_1683 NETTRAN_DUMMY_1684 MUX2_X1 
XU739 n724 n723 n458 n725 NETTRAN_DUMMY_1685 NETTRAN_DUMMY_1686 MUX2_X1 
XU738 n488 n513 n445 n724 NETTRAN_DUMMY_1687 NETTRAN_DUMMY_1688 MUX2_X1 
XU737 n535 n539 n445 n723 NETTRAN_DUMMY_1689 NETTRAN_DUMMY_1690 MUX2_X1 
XU736 n721 n718 n455 n722 NETTRAN_DUMMY_1691 NETTRAN_DUMMY_1692 MUX2_X1 
XU735 n720 n719 n458 n721 NETTRAN_DUMMY_1693 NETTRAN_DUMMY_1694 MUX2_X1 
XU734 n569 n536 n445 n720 NETTRAN_DUMMY_1695 NETTRAN_DUMMY_1696 MUX2_X1 
XU733 n480 n513 n445 n719 NETTRAN_DUMMY_1697 NETTRAN_DUMMY_1698 MUX2_X1 
XU732 n717 n716 n458 n718 NETTRAN_DUMMY_1699 NETTRAN_DUMMY_1700 MUX2_X1 
XU730 n531 n516 n445 n716 NETTRAN_DUMMY_1701 NETTRAN_DUMMY_1702 MUX2_X1 
XU729 n713 n714 n497 n715 NETTRAN_DUMMY_1703 NETTRAN_DUMMY_1704 MUX2_X1 
XU727 n711 n712 n452 n713 NETTRAN_DUMMY_1705 NETTRAN_DUMMY_1706 MUX2_X1 
XU725 n710 n709 n468 n711 NETTRAN_DUMMY_1707 NETTRAN_DUMMY_1708 MUX2_X1 
XU939 n923 n922 n477 n924 NETTRAN_DUMMY_1709 NETTRAN_DUMMY_1710 MUX2_X1 
XU938 n554 n1545 n500 n923 NETTRAN_DUMMY_1711 NETTRAN_DUMMY_1712 MUX2_X1 
XU937 n548 n1818 n500 n922 NETTRAN_DUMMY_1713 NETTRAN_DUMMY_1714 MUX2_X1 
XU936 n920 n913 n439 n921 NETTRAN_DUMMY_1715 NETTRAN_DUMMY_1716 MUX2_X1 
XU935 n919 n916 n454 n920 NETTRAN_DUMMY_1717 NETTRAN_DUMMY_1718 MUX2_X1 
XU934 n918 n917 n477 n919 NETTRAN_DUMMY_1719 NETTRAN_DUMMY_1720 MUX2_X1 
XU933 n563 n760 n507 n918 NETTRAN_DUMMY_1721 NETTRAN_DUMMY_1722 MUX2_X1 
XU932 n1796 n1815 n499 n917 NETTRAN_DUMMY_1723 NETTRAN_DUMMY_1724 MUX2_X1 
XU931 n915 n914 n475 n916 NETTRAN_DUMMY_1725 NETTRAN_DUMMY_1726 MUX2_X1 
XU930 n1853 n1767 n507 n915 NETTRAN_DUMMY_1727 NETTRAN_DUMMY_1728 MUX2_X1 
XU929 n1520 n548 n507 n914 NETTRAN_DUMMY_1729 NETTRAN_DUMMY_1730 MUX2_X1 
XU928 n911 n912 n454 n913 NETTRAN_DUMMY_1731 NETTRAN_DUMMY_1732 MUX2_X1 
XU926 n910 n909 n477 n911 NETTRAN_DUMMY_1733 NETTRAN_DUMMY_1734 MUX2_X1 
XU924 n1779 n608 n507 n909 NETTRAN_DUMMY_1735 NETTRAN_DUMMY_1736 MUX2_X1 
XU923 n1542 n523 n499 n908 NETTRAN_DUMMY_1737 NETTRAN_DUMMY_1738 MUX2_X1 
XU922 n907 n892 n433 d[20] NETTRAN_DUMMY_1739 NETTRAN_DUMMY_1740 MUX2_X1 
XU921 n906 n900 n443 n907 NETTRAN_DUMMY_1741 NETTRAN_DUMMY_1742 MUX2_X1 
XU920 n905 n902 n454 n906 NETTRAN_DUMMY_1743 NETTRAN_DUMMY_1744 MUX2_X1 
XU919 n904 n903 n475 n905 NETTRAN_DUMMY_1745 NETTRAN_DUMMY_1746 MUX2_X1 
XU918 n1775 n556 n507 n904 NETTRAN_DUMMY_1747 NETTRAN_DUMMY_1748 MUX2_X1 
XU917 n1785 n1745 n507 n903 NETTRAN_DUMMY_1749 NETTRAN_DUMMY_1750 MUX2_X1 
XU916 n901 n555 n477 n902 NETTRAN_DUMMY_1751 NETTRAN_DUMMY_1752 MUX2_X1 
XU915 n557 n488 n499 n901 NETTRAN_DUMMY_1753 NETTRAN_DUMMY_1754 MUX2_X1 
XU914 n899 n895 n454 n900 NETTRAN_DUMMY_1755 NETTRAN_DUMMY_1756 MUX2_X1 
XU913 n898 n896 n475 n899 NETTRAN_DUMMY_1757 NETTRAN_DUMMY_1758 MUX2_X1 
XU912 n517 n897 n507 n898 NETTRAN_DUMMY_1759 NETTRAN_DUMMY_1760 MUX2_X1 
XU910 n562 n591 n507 n896 NETTRAN_DUMMY_1761 NETTRAN_DUMMY_1762 MUX2_X1 
XU909 n894 n893 n475 n895 NETTRAN_DUMMY_1763 NETTRAN_DUMMY_1764 MUX2_X1 
XU908 n1522 n603 n507 n894 NETTRAN_DUMMY_1765 NETTRAN_DUMMY_1766 MUX2_X1 
XU907 n1789 n1784 n507 n893 NETTRAN_DUMMY_1767 NETTRAN_DUMMY_1768 MUX2_X1 
XU906 n891 n885 n445 n892 NETTRAN_DUMMY_1769 NETTRAN_DUMMY_1770 MUX2_X1 
XU905 n890 n888 n455 n891 NETTRAN_DUMMY_1771 NETTRAN_DUMMY_1772 MUX2_X1 
XU904 n512 n889 n475 n890 NETTRAN_DUMMY_1773 NETTRAN_DUMMY_1774 MUX2_X1 
XU903 n1333 n523 n507 n889 NETTRAN_DUMMY_1775 NETTRAN_DUMMY_1776 MUX2_X1 
XU902 n887 n886 n475 n888 NETTRAN_DUMMY_1777 NETTRAN_DUMMY_1778 MUX2_X1 
XU901 n563 n542 n507 n887 NETTRAN_DUMMY_1779 NETTRAN_DUMMY_1780 MUX2_X1 
XU900 n1741 n1831 n507 n886 NETTRAN_DUMMY_1781 NETTRAN_DUMMY_1782 MUX2_X1 
XU899 n882 n883 n448 n885 NETTRAN_DUMMY_1783 NETTRAN_DUMMY_1784 MUX2_X1 
XU897 n881 n880 n473 n882 NETTRAN_DUMMY_1785 NETTRAN_DUMMY_1786 MUX2_X1 
XU896 n526 n520 n497 n881 NETTRAN_DUMMY_1787 NETTRAN_DUMMY_1788 MUX2_X1 
XU895 n527 n538 n507 n880 NETTRAN_DUMMY_1789 NETTRAN_DUMMY_1790 MUX2_X1 
XU894 n879 n864 n433 d[1] NETTRAN_DUMMY_1791 NETTRAN_DUMMY_1792 MUX2_X1 
XU893 n878 n871 n439 n879 NETTRAN_DUMMY_1793 NETTRAN_DUMMY_1794 MUX2_X1 
XU892 n877 n874 n452 n878 NETTRAN_DUMMY_1795 NETTRAN_DUMMY_1796 MUX2_X1 
XU891 n876 n875 n499 n877 NETTRAN_DUMMY_1797 NETTRAN_DUMMY_1798 MUX2_X1 
XU890 n1815 n1674 n475 n876 NETTRAN_DUMMY_1799 NETTRAN_DUMMY_1800 MUX2_X1 
XU889 n1761 n1767 n475 n875 NETTRAN_DUMMY_1801 NETTRAN_DUMMY_1802 MUX2_X1 
XU888 n872 n873 n503 n874 NETTRAN_DUMMY_1803 NETTRAN_DUMMY_1804 MUX2_X1 
XU886 n547 n1759 n473 n872 NETTRAN_DUMMY_1805 NETTRAN_DUMMY_1806 MUX2_X1 
XU885 n870 n867 n452 n871 NETTRAN_DUMMY_1807 NETTRAN_DUMMY_1808 MUX2_X1 
XU884 n869 n868 n503 n870 NETTRAN_DUMMY_1809 NETTRAN_DUMMY_1810 MUX2_X1 
XU882 n525 n1853 n475 n868 NETTRAN_DUMMY_1811 NETTRAN_DUMMY_1812 MUX2_X1 
XU881 n866 n865 n503 n867 NETTRAN_DUMMY_1813 NETTRAN_DUMMY_1814 MUX2_X1 
XU880 n1759 n1541 n473 n866 NETTRAN_DUMMY_1815 NETTRAN_DUMMY_1816 MUX2_X1 
XU879 n1520 n581 n473 n865 NETTRAN_DUMMY_1817 NETTRAN_DUMMY_1818 MUX2_X1 
XU878 n863 n856 n439 n864 NETTRAN_DUMMY_1819 NETTRAN_DUMMY_1820 MUX2_X1 
XU877 n862 n859 n452 n863 NETTRAN_DUMMY_1821 NETTRAN_DUMMY_1822 MUX2_X1 
XU876 n861 n860 n503 n862 NETTRAN_DUMMY_1823 NETTRAN_DUMMY_1824 MUX2_X1 
XU875 n575 n557 n462 n861 NETTRAN_DUMMY_1825 NETTRAN_DUMMY_1826 MUX2_X1 
XU874 n1778 n1535 n473 n860 NETTRAN_DUMMY_1827 NETTRAN_DUMMY_1828 MUX2_X1 
XU873 n858 n857 n503 n859 NETTRAN_DUMMY_1829 NETTRAN_DUMMY_1830 MUX2_X1 
XU872 n515 n410 n462 n858 NETTRAN_DUMMY_1831 NETTRAN_DUMMY_1832 MUX2_X1 
XU871 n1779 n760 n475 n857 NETTRAN_DUMMY_1833 NETTRAN_DUMMY_1834 MUX2_X1 
XU870 n853 n854 n452 n856 NETTRAN_DUMMY_1835 NETTRAN_DUMMY_1836 MUX2_X1 
XU868 n852 n851 n507 n853 NETTRAN_DUMMY_1837 NETTRAN_DUMMY_1838 MUX2_X1 
XU867 n1525 n1533 n475 n852 NETTRAN_DUMMY_1839 NETTRAN_DUMMY_1840 MUX2_X1 
XU866 n1674 n1501 n475 n851 NETTRAN_DUMMY_1841 NETTRAN_DUMMY_1842 MUX2_X1 
XU865 n850 n834 n433 d[19] NETTRAN_DUMMY_1843 NETTRAN_DUMMY_1844 MUX2_X1 
XU864 n849 n842 n455 n850 NETTRAN_DUMMY_1845 NETTRAN_DUMMY_1846 MUX2_X1 
XU863 n848 n845 n495 n849 NETTRAN_DUMMY_1847 NETTRAN_DUMMY_1848 MUX2_X1 
XU862 n847 n846 n458 n848 NETTRAN_DUMMY_1849 NETTRAN_DUMMY_1850 MUX2_X1 
XU861 n1533 n1521 n443 n847 NETTRAN_DUMMY_1851 NETTRAN_DUMMY_1852 MUX2_X1 
XU860 n529 n1776 n443 n846 NETTRAN_DUMMY_1853 NETTRAN_DUMMY_1854 MUX2_X1 
XU859 n843 n844 n458 n845 NETTRAN_DUMMY_1855 NETTRAN_DUMMY_1856 MUX2_X1 
XU857 n1801 n1817 n443 n843 NETTRAN_DUMMY_1857 NETTRAN_DUMMY_1858 MUX2_X1 
XU856 n841 n838 n495 n842 NETTRAN_DUMMY_1859 NETTRAN_DUMMY_1860 MUX2_X1 
XU855 n840 n839 n458 n841 NETTRAN_DUMMY_1861 NETTRAN_DUMMY_1862 MUX2_X1 
XU854 n1523 n573 n443 n840 NETTRAN_DUMMY_1863 NETTRAN_DUMMY_1864 MUX2_X1 
XU853 n492 n1530 n445 n839 NETTRAN_DUMMY_1865 NETTRAN_DUMMY_1866 MUX2_X1 
XU852 n835 n836 n458 n838 NETTRAN_DUMMY_1867 NETTRAN_DUMMY_1868 MUX2_X1 
XU850 n1545 n1523 n443 n835 NETTRAN_DUMMY_1869 NETTRAN_DUMMY_1870 MUX2_X1 
XU849 n833 n826 n455 n834 NETTRAN_DUMMY_1871 NETTRAN_DUMMY_1872 MUX2_X1 
XU848 n832 n829 n495 n833 NETTRAN_DUMMY_1873 NETTRAN_DUMMY_1874 MUX2_X1 
XU847 n831 n830 n471 n832 NETTRAN_DUMMY_1875 NETTRAN_DUMMY_1876 MUX2_X1 
XU846 n1754 n1500 n443 n831 NETTRAN_DUMMY_1877 NETTRAN_DUMMY_1878 MUX2_X1 
XU845 n1850 n1814 n443 n830 NETTRAN_DUMMY_1879 NETTRAN_DUMMY_1880 MUX2_X1 
XU844 n828 n827 n471 n829 NETTRAN_DUMMY_1881 NETTRAN_DUMMY_1882 MUX2_X1 
XU843 n1817 n531 n443 n828 NETTRAN_DUMMY_1883 NETTRAN_DUMMY_1884 MUX2_X1 
XU842 n1808 n1776 n443 n827 NETTRAN_DUMMY_1885 NETTRAN_DUMMY_1886 MUX2_X1 
XU841 n824 n825 n495 n826 NETTRAN_DUMMY_1887 NETTRAN_DUMMY_1888 MUX2_X1 
XU839 n822 n823 n458 n824 NETTRAN_DUMMY_1889 NETTRAN_DUMMY_1890 MUX2_X1 
XU837 n1772 n1781 n443 n822 NETTRAN_DUMMY_1891 NETTRAN_DUMMY_1892 MUX2_X1 
XU836 n601 n629 n443 n821 NETTRAN_DUMMY_1893 NETTRAN_DUMMY_1894 MUX2_X1 
XU1039 n1020 n1017 n503 n1021 NETTRAN_DUMMY_1895 NETTRAN_DUMMY_1896 MUX2_X1 
XU1038 n1019 n1018 n462 n1020 NETTRAN_DUMMY_1897 NETTRAN_DUMMY_1898 MUX2_X1 
XU1037 n555 n515 n435 n1019 NETTRAN_DUMMY_1899 NETTRAN_DUMMY_1900 MUX2_X1 
XU1036 n615 n1768 n435 n1018 NETTRAN_DUMMY_1901 NETTRAN_DUMMY_1902 MUX2_X1 
XU1035 n1016 n1015 n462 n1017 NETTRAN_DUMMY_1903 NETTRAN_DUMMY_1904 MUX2_X1 
XU1034 n897 n1544 n435 n1016 NETTRAN_DUMMY_1905 NETTRAN_DUMMY_1906 MUX2_X1 
XU1033 n564 n1746 n435 n1015 NETTRAN_DUMMY_1907 NETTRAN_DUMMY_1908 MUX2_X1 
XU1032 n1013 n1010 n503 n1014 NETTRAN_DUMMY_1909 NETTRAN_DUMMY_1910 MUX2_X1 
XU1031 n1012 n1011 n464 n1013 NETTRAN_DUMMY_1911 NETTRAN_DUMMY_1912 MUX2_X1 
XU1030 n1752 n1747 n435 n1012 NETTRAN_DUMMY_1913 NETTRAN_DUMMY_1914 MUX2_X1 
XU1029 n1352 n562 n435 n1011 NETTRAN_DUMMY_1915 NETTRAN_DUMMY_1916 MUX2_X1 
XU1028 n1009 n1008 n462 n1010 NETTRAN_DUMMY_1917 NETTRAN_DUMMY_1918 MUX2_X1 
XU1027 n593 n617 n435 n1009 NETTRAN_DUMMY_1919 NETTRAN_DUMMY_1920 MUX2_X1 
XU1026 n537 n493 n435 n1008 NETTRAN_DUMMY_1921 NETTRAN_DUMMY_1922 MUX2_X1 
XU1025 n1006 n999 n452 n1007 NETTRAN_DUMMY_1923 NETTRAN_DUMMY_1924 MUX2_X1 
XU1024 n1005 n1002 n507 n1006 NETTRAN_DUMMY_1925 NETTRAN_DUMMY_1926 MUX2_X1 
XU1023 n1004 n1003 n475 n1005 NETTRAN_DUMMY_1927 NETTRAN_DUMMY_1928 MUX2_X1 
XU1022 n1756 n584 n435 n1004 NETTRAN_DUMMY_1929 NETTRAN_DUMMY_1930 MUX2_X1 
XU1021 n566 n629 n435 n1003 NETTRAN_DUMMY_1931 NETTRAN_DUMMY_1932 MUX2_X1 
XU1020 n1001 n1000 n475 n1002 NETTRAN_DUMMY_1933 NETTRAN_DUMMY_1934 MUX2_X1 
XU1019 n1840 n1745 n435 n1001 NETTRAN_DUMMY_1935 NETTRAN_DUMMY_1936 MUX2_X1 
XU1018 n579 n609 n435 n1000 NETTRAN_DUMMY_1937 NETTRAN_DUMMY_1938 MUX2_X1 
XU1017 n998 n995 n503 n999 NETTRAN_DUMMY_1939 NETTRAN_DUMMY_1940 MUX2_X1 
XU1016 n996 n997 n462 n998 NETTRAN_DUMMY_1941 NETTRAN_DUMMY_1942 MUX2_X1 
XU1014 n1755 n615 n435 n996 NETTRAN_DUMMY_1943 NETTRAN_DUMMY_1944 MUX2_X1 
XU1013 n994 n993 n473 n995 NETTRAN_DUMMY_1945 NETTRAN_DUMMY_1946 MUX2_X1 
XU1010 n992 n977 n435 d[23] NETTRAN_DUMMY_1947 NETTRAN_DUMMY_1948 MUX2_X1 
XU1009 n991 n984 n439 n992 NETTRAN_DUMMY_1949 NETTRAN_DUMMY_1950 MUX2_X1 
XU1008 n990 n987 n454 n991 NETTRAN_DUMMY_1951 NETTRAN_DUMMY_1952 MUX2_X1 
XU1007 n989 n988 n499 n990 NETTRAN_DUMMY_1953 NETTRAN_DUMMY_1954 MUX2_X1 
XU1006 n1529 n572 n477 n989 NETTRAN_DUMMY_1955 NETTRAN_DUMMY_1956 MUX2_X1 
XU1005 n1777 n612 n477 n988 NETTRAN_DUMMY_1957 NETTRAN_DUMMY_1958 MUX2_X1 
XU1004 n986 n985 n499 n987 NETTRAN_DUMMY_1959 NETTRAN_DUMMY_1960 MUX2_X1 
XU1003 n571 n1775 n477 n986 NETTRAN_DUMMY_1961 NETTRAN_DUMMY_1962 MUX2_X1 
XU1002 n1529 n606 n477 n985 NETTRAN_DUMMY_1963 NETTRAN_DUMMY_1964 MUX2_X1 
XU1001 n983 n980 n454 n984 NETTRAN_DUMMY_1965 NETTRAN_DUMMY_1966 MUX2_X1 
XU1000 n982 n981 n499 n983 NETTRAN_DUMMY_1967 NETTRAN_DUMMY_1968 MUX2_X1 
XU999 n492 n586 n477 n982 NETTRAN_DUMMY_1969 NETTRAN_DUMMY_1970 MUX2_X1 
XU998 n571 n583 n477 n981 NETTRAN_DUMMY_1971 NETTRAN_DUMMY_1972 MUX2_X1 
XU997 n979 n978 n499 n980 NETTRAN_DUMMY_1973 NETTRAN_DUMMY_1974 MUX2_X1 
XU996 n1780 n565 n462 n979 NETTRAN_DUMMY_1975 NETTRAN_DUMMY_1976 MUX2_X1 
XU995 n1783 n602 n462 n978 NETTRAN_DUMMY_1977 NETTRAN_DUMMY_1978 MUX2_X1 
XU994 n976 n970 n439 n977 NETTRAN_DUMMY_1979 NETTRAN_DUMMY_1980 MUX2_X1 
XU993 n975 n973 n452 n976 NETTRAN_DUMMY_1981 NETTRAN_DUMMY_1982 MUX2_X1 
XU992 n547 n974 n428 n975 NETTRAN_DUMMY_1983 NETTRAN_DUMMY_1984 MUX2_X1 
XU991 n544 n1754 n507 n974 NETTRAN_DUMMY_1985 NETTRAN_DUMMY_1986 MUX2_X1 
XU990 n972 n971 n507 n973 NETTRAN_DUMMY_1987 NETTRAN_DUMMY_1988 MUX2_X1 
XU989 n530 n1797 n475 n972 NETTRAN_DUMMY_1989 NETTRAN_DUMMY_1990 MUX2_X1 
XU988 n1521 n520 n475 n971 NETTRAN_DUMMY_1991 NETTRAN_DUMMY_1992 MUX2_X1 
XU987 n968 n969 n452 n970 NETTRAN_DUMMY_1993 NETTRAN_DUMMY_1994 MUX2_X1 
XU985 n967 n966 n503 n968 NETTRAN_DUMMY_1995 NETTRAN_DUMMY_1996 MUX2_X1 
XU983 n591 n1754 n473 n966 NETTRAN_DUMMY_1997 NETTRAN_DUMMY_1998 MUX2_X1 
XU982 n1812 n492 n507 n965 NETTRAN_DUMMY_1999 NETTRAN_DUMMY_2000 MUX2_X1 
XU981 n964 n949 n435 d[22] NETTRAN_DUMMY_2001 NETTRAN_DUMMY_2002 MUX2_X1 
XU980 n963 n956 n439 n964 NETTRAN_DUMMY_2003 NETTRAN_DUMMY_2004 MUX2_X1 
XU979 n962 n959 n452 n963 NETTRAN_DUMMY_2005 NETTRAN_DUMMY_2006 MUX2_X1 
XU978 n961 n960 n507 n962 NETTRAN_DUMMY_2007 NETTRAN_DUMMY_2008 MUX2_X1 
XU977 n526 n516 n473 n961 NETTRAN_DUMMY_2009 NETTRAN_DUMMY_2010 MUX2_X1 
XU976 n522 n1743 n475 n960 NETTRAN_DUMMY_2011 NETTRAN_DUMMY_2012 MUX2_X1 
XU975 n958 n957 n507 n959 NETTRAN_DUMMY_2013 NETTRAN_DUMMY_2014 MUX2_X1 
XU974 n1799 n1790 n475 n958 NETTRAN_DUMMY_2015 NETTRAN_DUMMY_2016 MUX2_X1 
XU973 n1541 n595 n475 n957 NETTRAN_DUMMY_2017 NETTRAN_DUMMY_2018 MUX2_X1 
XU972 n955 n952 n454 n956 NETTRAN_DUMMY_2019 NETTRAN_DUMMY_2020 MUX2_X1 
XU971 n954 n953 n499 n955 NETTRAN_DUMMY_2021 NETTRAN_DUMMY_2022 MUX2_X1 
XU970 n1845 n1759 n477 n954 NETTRAN_DUMMY_2023 NETTRAN_DUMMY_2024 MUX2_X1 
XU969 n1318 n565 n462 n953 NETTRAN_DUMMY_2025 NETTRAN_DUMMY_2026 MUX2_X1 
XU968 n951 n950 n499 n952 NETTRAN_DUMMY_2027 NETTRAN_DUMMY_2028 MUX2_X1 
XU967 n1825 n1762 n477 n951 NETTRAN_DUMMY_2029 NETTRAN_DUMMY_2030 MUX2_X1 
XU966 n527 n588 n477 n950 NETTRAN_DUMMY_2031 NETTRAN_DUMMY_2032 MUX2_X1 
XU965 n948 n941 n439 n949 NETTRAN_DUMMY_2033 NETTRAN_DUMMY_2034 MUX2_X1 
XU964 n947 n944 n454 n948 NETTRAN_DUMMY_2035 NETTRAN_DUMMY_2036 MUX2_X1 
XU963 n946 n945 n499 n947 NETTRAN_DUMMY_2037 NETTRAN_DUMMY_2038 MUX2_X1 
XU962 n570 n1500 n462 n946 NETTRAN_DUMMY_2039 NETTRAN_DUMMY_2040 MUX2_X1 
XU961 n776 n564 n462 n945 NETTRAN_DUMMY_2041 NETTRAN_DUMMY_2042 MUX2_X1 
XU960 n943 n942 n499 n944 NETTRAN_DUMMY_2043 NETTRAN_DUMMY_2044 MUX2_X1 
XU959 n608 n573 n477 n943 NETTRAN_DUMMY_2045 NETTRAN_DUMMY_2046 MUX2_X1 
XU958 n1808 n542 n477 n942 NETTRAN_DUMMY_2047 NETTRAN_DUMMY_2048 MUX2_X1 
XU957 n939 n940 n454 n941 NETTRAN_DUMMY_2049 NETTRAN_DUMMY_2050 MUX2_X1 
XU955 n938 n937 n499 n939 NETTRAN_DUMMY_2051 NETTRAN_DUMMY_2052 MUX2_X1 
XU954 n555 n601 n477 n938 NETTRAN_DUMMY_2053 NETTRAN_DUMMY_2054 MUX2_X1 
XU953 n583 n1787 n477 n937 NETTRAN_DUMMY_2055 NETTRAN_DUMMY_2056 MUX2_X1 
XU952 n602 n1526 n499 n936 NETTRAN_DUMMY_2057 NETTRAN_DUMMY_2058 MUX2_X1 
XU951 n935 n921 n435 d[21] NETTRAN_DUMMY_2059 NETTRAN_DUMMY_2060 MUX2_X1 
XU950 n934 n928 n443 n935 NETTRAN_DUMMY_2061 NETTRAN_DUMMY_2062 MUX2_X1 
XU949 n933 n930 n452 n934 NETTRAN_DUMMY_2063 NETTRAN_DUMMY_2064 MUX2_X1 
XU948 n932 n931 n475 n933 NETTRAN_DUMMY_2065 NETTRAN_DUMMY_2066 MUX2_X1 
XU946 n562 n550 n507 n931 NETTRAN_DUMMY_2067 NETTRAN_DUMMY_2068 MUX2_X1 
XU945 n929 n1806 n475 n930 NETTRAN_DUMMY_2069 NETTRAN_DUMMY_2070 MUX2_X1 
XU944 n1760 n583 n507 n929 NETTRAN_DUMMY_2071 NETTRAN_DUMMY_2072 MUX2_X1 
XU943 n927 n924 n454 n928 NETTRAN_DUMMY_2073 NETTRAN_DUMMY_2074 MUX2_X1 
XU942 n926 n925 n477 n927 NETTRAN_DUMMY_2075 NETTRAN_DUMMY_2076 MUX2_X1 
XU941 n410 n517 n499 n926 NETTRAN_DUMMY_2077 NETTRAN_DUMMY_2078 MUX2_X1 
XU940 n1532 n593 n500 n925 NETTRAN_DUMMY_2079 NETTRAN_DUMMY_2080 MUX2_X1 
XU1142 n523 n567 n462 n1124 NETTRAN_DUMMY_2081 NETTRAN_DUMMY_2082 MUX2_X1 
XU1141 n1122 n1119 n452 n1123 NETTRAN_DUMMY_2083 NETTRAN_DUMMY_2084 MUX2_X1 
XU1140 n1121 n1120 n503 n1122 NETTRAN_DUMMY_2085 NETTRAN_DUMMY_2086 MUX2_X1 
XU1139 n551 n1543 n473 n1121 NETTRAN_DUMMY_2087 NETTRAN_DUMMY_2088 MUX2_X1 
XU1138 n1538 n567 n462 n1120 NETTRAN_DUMMY_2089 NETTRAN_DUMMY_2090 MUX2_X1 
XU1137 n1118 n1667 n503 n1119 NETTRAN_DUMMY_2091 NETTRAN_DUMMY_2092 MUX2_X1 
XU1136 n539 n1826 n462 n1118 NETTRAN_DUMMY_2093 NETTRAN_DUMMY_2094 MUX2_X1 
XU1135 n1114 n1115 n439 n1117 NETTRAN_DUMMY_2095 NETTRAN_DUMMY_2096 MUX2_X1 
XU1133 n1113 n1111 n452 n1114 NETTRAN_DUMMY_2097 NETTRAN_DUMMY_2098 MUX2_X1 
XU1132 n1112 n623 n503 n1113 NETTRAN_DUMMY_2099 NETTRAN_DUMMY_2100 MUX2_X1 
XU1130 n1110 n513 n503 n1111 NETTRAN_DUMMY_2101 NETTRAN_DUMMY_2102 MUX2_X1 
XU1128 n623 n1521 n452 n1109 NETTRAN_DUMMY_2103 NETTRAN_DUMMY_2104 MUX2_X1 
XU1127 n501 n624 n452 n1108 NETTRAN_DUMMY_2105 NETTRAN_DUMMY_2106 MUX2_X1 
XU1126 n1107 n1092 n435 d[27] NETTRAN_DUMMY_2107 NETTRAN_DUMMY_2108 MUX2_X1 
XU1125 n1106 n1099 n439 n1107 NETTRAN_DUMMY_2109 NETTRAN_DUMMY_2110 MUX2_X1 
XU1124 n1105 n1102 n453 n1106 NETTRAN_DUMMY_2111 NETTRAN_DUMMY_2112 MUX2_X1 
XU1123 n1104 n1103 n500 n1105 NETTRAN_DUMMY_2113 NETTRAN_DUMMY_2114 MUX2_X1 
XU1122 n1749 n1825 n464 n1104 NETTRAN_DUMMY_2115 NETTRAN_DUMMY_2116 MUX2_X1 
XU1121 n565 n545 n464 n1103 NETTRAN_DUMMY_2117 NETTRAN_DUMMY_2118 MUX2_X1 
XU1120 n1101 n1100 n500 n1102 NETTRAN_DUMMY_2119 NETTRAN_DUMMY_2120 MUX2_X1 
XU1119 n548 n620 n464 n1101 NETTRAN_DUMMY_2121 NETTRAN_DUMMY_2122 MUX2_X1 
XU1118 n1841 n1759 n464 n1100 NETTRAN_DUMMY_2123 NETTRAN_DUMMY_2124 MUX2_X1 
XU1117 n1098 n1095 n452 n1099 NETTRAN_DUMMY_2125 NETTRAN_DUMMY_2126 MUX2_X1 
XU1116 n1097 n1096 n503 n1098 NETTRAN_DUMMY_2127 NETTRAN_DUMMY_2128 MUX2_X1 
XU1115 n598 n557 n462 n1097 NETTRAN_DUMMY_2129 NETTRAN_DUMMY_2130 MUX2_X1 
XU1114 n410 n1805 n462 n1096 NETTRAN_DUMMY_2131 NETTRAN_DUMMY_2132 MUX2_X1 
XU1113 n1093 n1094 n503 n1095 NETTRAN_DUMMY_2133 NETTRAN_DUMMY_2134 MUX2_X1 
XU1111 n410 n1826 n462 n1093 NETTRAN_DUMMY_2135 NETTRAN_DUMMY_2136 MUX2_X1 
XU1110 n1091 n1085 n439 n1092 NETTRAN_DUMMY_2137 NETTRAN_DUMMY_2138 MUX2_X1 
XU1109 n1090 n1087 n454 n1091 NETTRAN_DUMMY_2139 NETTRAN_DUMMY_2140 MUX2_X1 
XU1108 n1089 n1088 n499 n1090 NETTRAN_DUMMY_2141 NETTRAN_DUMMY_2142 MUX2_X1 
XU1107 n1808 n536 n462 n1089 NETTRAN_DUMMY_2143 NETTRAN_DUMMY_2144 MUX2_X1 
XU1106 n1542 n581 n462 n1088 NETTRAN_DUMMY_2145 NETTRAN_DUMMY_2146 MUX2_X1 
XU1105 n1538 n1086 n428 n1087 NETTRAN_DUMMY_2147 NETTRAN_DUMMY_2148 MUX2_X1 
XU1103 n1082 n1083 n454 n1085 NETTRAN_DUMMY_2149 NETTRAN_DUMMY_2150 MUX2_X1 
XU1101 n1081 n1080 n499 n1082 NETTRAN_DUMMY_2151 NETTRAN_DUMMY_2152 MUX2_X1 
XU1100 n515 n612 n462 n1081 NETTRAN_DUMMY_2153 NETTRAN_DUMMY_2154 MUX2_X1 
XU1099 n593 n581 n462 n1080 NETTRAN_DUMMY_2155 NETTRAN_DUMMY_2156 MUX2_X1 
XU1098 n1079 n1064 n435 d[26] NETTRAN_DUMMY_2157 NETTRAN_DUMMY_2158 MUX2_X1 
XU1097 n1078 n1071 n439 n1079 NETTRAN_DUMMY_2159 NETTRAN_DUMMY_2160 MUX2_X1 
XU1096 n1077 n1074 n454 n1078 NETTRAN_DUMMY_2161 NETTRAN_DUMMY_2162 MUX2_X1 
XU1095 n1076 n1075 n500 n1077 NETTRAN_DUMMY_2163 NETTRAN_DUMMY_2164 MUX2_X1 
XU1094 n1771 n523 n464 n1076 NETTRAN_DUMMY_2165 NETTRAN_DUMMY_2166 MUX2_X1 
XU1093 n599 n1333 n464 n1075 NETTRAN_DUMMY_2167 NETTRAN_DUMMY_2168 MUX2_X1 
XU1092 n1073 n1072 n499 n1074 NETTRAN_DUMMY_2169 NETTRAN_DUMMY_2170 MUX2_X1 
XU1091 n596 n560 n477 n1073 NETTRAN_DUMMY_2171 NETTRAN_DUMMY_2172 MUX2_X1 
XU1090 n1742 n1779 n475 n1072 NETTRAN_DUMMY_2173 NETTRAN_DUMMY_2174 MUX2_X1 
XU1089 n1069 n1067 n454 n1071 NETTRAN_DUMMY_2175 NETTRAN_DUMMY_2176 MUX2_X1 
XU1088 n1068 n1070 n499 n1069 NETTRAN_DUMMY_2177 NETTRAN_DUMMY_2178 MUX2_X1 
XU1087 n602 n629 n462 n1068 NETTRAN_DUMMY_2179 NETTRAN_DUMMY_2180 MUX2_X1 
XU1086 n1066 n1065 n499 n1067 NETTRAN_DUMMY_2181 NETTRAN_DUMMY_2182 MUX2_X1 
XU1085 n1846 n523 n462 n1066 NETTRAN_DUMMY_2183 NETTRAN_DUMMY_2184 MUX2_X1 
XU1084 n1748 n619 n462 n1065 NETTRAN_DUMMY_2185 NETTRAN_DUMMY_2186 MUX2_X1 
XU1083 n1063 n1056 n439 n1064 NETTRAN_DUMMY_2187 NETTRAN_DUMMY_2188 MUX2_X1 
XU1082 n1062 n1059 n452 n1063 NETTRAN_DUMMY_2189 NETTRAN_DUMMY_2190 MUX2_X1 
XU1081 n1061 n1060 n503 n1062 NETTRAN_DUMMY_2191 NETTRAN_DUMMY_2192 MUX2_X1 
XU1079 n1776 n567 n462 n1060 NETTRAN_DUMMY_2193 NETTRAN_DUMMY_2194 MUX2_X1 
XU1078 n1058 n1057 n499 n1059 NETTRAN_DUMMY_2195 NETTRAN_DUMMY_2196 MUX2_X1 
XU1077 n566 n1827 n462 n1058 NETTRAN_DUMMY_2197 NETTRAN_DUMMY_2198 MUX2_X1 
XU1076 n1538 n1541 n462 n1057 NETTRAN_DUMMY_2199 NETTRAN_DUMMY_2200 MUX2_X1 
XU1075 n1054 n1055 n454 n1056 NETTRAN_DUMMY_2201 NETTRAN_DUMMY_2202 MUX2_X1 
XU1073 n1053 n1052 n499 n1054 NETTRAN_DUMMY_2203 NETTRAN_DUMMY_2204 MUX2_X1 
XU1072 IN1 n601 n462 n1053 NETTRAN_DUMMY_2205 NETTRAN_DUMMY_2206 MUX2_X1 
XU1071 n612 n1833 n462 n1052 NETTRAN_DUMMY_2207 NETTRAN_DUMMY_2208 MUX2_X1 
XU1070 n536 n628 n499 n1051 NETTRAN_DUMMY_2209 NETTRAN_DUMMY_2210 MUX2_X1 
XU1069 n1050 n1035 n435 d[25] NETTRAN_DUMMY_2211 NETTRAN_DUMMY_2212 MUX2_X1 
XU1068 n1049 n1042 n439 n1050 NETTRAN_DUMMY_2213 NETTRAN_DUMMY_2214 MUX2_X1 
XU1067 n1048 n1045 n452 n1049 NETTRAN_DUMMY_2215 NETTRAN_DUMMY_2216 MUX2_X1 
XU1066 n1047 n1046 n503 n1048 NETTRAN_DUMMY_2217 NETTRAN_DUMMY_2218 MUX2_X1 
XU1065 n535 n567 n462 n1047 NETTRAN_DUMMY_2219 NETTRAN_DUMMY_2220 MUX2_X1 
XU1064 n592 n897 n473 n1046 NETTRAN_DUMMY_2221 NETTRAN_DUMMY_2222 MUX2_X1 
XU1063 n1044 n1043 n503 n1045 NETTRAN_DUMMY_2223 NETTRAN_DUMMY_2224 MUX2_X1 
XU1062 n1826 n566 n462 n1044 NETTRAN_DUMMY_2225 NETTRAN_DUMMY_2226 MUX2_X1 
XU1061 n1805 n598 n462 n1043 NETTRAN_DUMMY_2227 NETTRAN_DUMMY_2228 MUX2_X1 
XU1060 n1041 n1038 n453 n1042 NETTRAN_DUMMY_2229 NETTRAN_DUMMY_2230 MUX2_X1 
XU1059 n1040 n1039 n500 n1041 NETTRAN_DUMMY_2231 NETTRAN_DUMMY_2232 MUX2_X1 
XU1058 n1818 n1795 n475 n1040 NETTRAN_DUMMY_2233 NETTRAN_DUMMY_2234 MUX2_X1 
XU1057 n1333 n1824 n475 n1039 NETTRAN_DUMMY_2235 NETTRAN_DUMMY_2236 MUX2_X1 
XU1056 n1037 n1036 n500 n1038 NETTRAN_DUMMY_2237 NETTRAN_DUMMY_2238 MUX2_X1 
XU1055 n605 n1841 n464 n1037 NETTRAN_DUMMY_2239 NETTRAN_DUMMY_2240 MUX2_X1 
XU1054 n613 n576 n475 n1036 NETTRAN_DUMMY_2241 NETTRAN_DUMMY_2242 MUX2_X1 
XU1053 n1034 n1028 n439 n1035 NETTRAN_DUMMY_2243 NETTRAN_DUMMY_2244 MUX2_X1 
XU1052 n1033 n1031 n454 n1034 NETTRAN_DUMMY_2245 NETTRAN_DUMMY_2246 MUX2_X1 
XU1051 n1672 n1032 n507 n1033 NETTRAN_DUMMY_2247 NETTRAN_DUMMY_2248 MUX2_X1 
XU1050 n1839 n573 n475 n1032 NETTRAN_DUMMY_2249 NETTRAN_DUMMY_2250 MUX2_X1 
XU1049 n1030 n1029 n499 n1031 NETTRAN_DUMMY_2251 NETTRAN_DUMMY_2252 MUX2_X1 
XU1048 n561 n1789 n462 n1030 NETTRAN_DUMMY_2253 NETTRAN_DUMMY_2254 MUX2_X1 
XU1047 n557 n533 n462 n1029 NETTRAN_DUMMY_2255 NETTRAN_DUMMY_2256 MUX2_X1 
XU1046 n1025 n1026 n454 n1028 NETTRAN_DUMMY_2257 NETTRAN_DUMMY_2258 MUX2_X1 
XU1044 n1024 n1023 n499 n1025 NETTRAN_DUMMY_2259 NETTRAN_DUMMY_2260 MUX2_X1 
XU1042 n601 n1826 n477 n1023 NETTRAN_DUMMY_2261 NETTRAN_DUMMY_2262 MUX2_X1 
XU1041 n1022 n1007 n439 d[24] NETTRAN_DUMMY_2263 NETTRAN_DUMMY_2264 MUX2_X1 
XU1040 n1021 n1014 n452 n1022 NETTRAN_DUMMY_2265 NETTRAN_DUMMY_2266 MUX2_X1 
XU1248 n1757 n1225 n466 n1226 NETTRAN_DUMMY_2267 NETTRAN_DUMMY_2268 MUX2_X1 
XU1247 n1318 n614 n502 n1225 NETTRAN_DUMMY_2269 NETTRAN_DUMMY_2270 MUX2_X1 
XU1246 n1223 n1222 n466 n1224 NETTRAN_DUMMY_2271 NETTRAN_DUMMY_2272 MUX2_X1 
XU1245 n610 n1772 n502 n1223 NETTRAN_DUMMY_2273 NETTRAN_DUMMY_2274 MUX2_X1 
XU1244 n528 n570 n500 n1222 NETTRAN_DUMMY_2275 NETTRAN_DUMMY_2276 MUX2_X1 
XU1243 n1220 n1217 n453 n1221 NETTRAN_DUMMY_2277 NETTRAN_DUMMY_2278 MUX2_X1 
XU1242 n1219 n1218 n466 n1220 NETTRAN_DUMMY_2279 NETTRAN_DUMMY_2280 MUX2_X1 
XU1241 n1783 n1532 n502 n1219 NETTRAN_DUMMY_2281 NETTRAN_DUMMY_2282 MUX2_X1 
XU1240 n625 n1333 n502 n1218 NETTRAN_DUMMY_2283 NETTRAN_DUMMY_2284 MUX2_X1 
XU1239 n1216 n1215 n466 n1217 NETTRAN_DUMMY_2285 NETTRAN_DUMMY_2286 MUX2_X1 
XU1238 n1811 n1534 n507 n1216 NETTRAN_DUMMY_2287 NETTRAN_DUMMY_2288 MUX2_X1 
XU1237 n1791 n606 n502 n1215 NETTRAN_DUMMY_2289 NETTRAN_DUMMY_2290 MUX2_X1 
XU1236 n1213 n1206 n442 n1214 NETTRAN_DUMMY_2291 NETTRAN_DUMMY_2292 MUX2_X1 
XU1235 n1212 n1209 n453 n1213 NETTRAN_DUMMY_2293 NETTRAN_DUMMY_2294 MUX2_X1 
XU1234 n1211 n1210 n466 n1212 NETTRAN_DUMMY_2295 NETTRAN_DUMMY_2296 MUX2_X1 
XU1233 n610 n615 n502 n1211 NETTRAN_DUMMY_2297 NETTRAN_DUMMY_2298 MUX2_X1 
XU1232 n1828 n1500 n502 n1210 NETTRAN_DUMMY_2299 NETTRAN_DUMMY_2300 MUX2_X1 
XU1231 n1208 n1207 n466 n1209 NETTRAN_DUMMY_2301 NETTRAN_DUMMY_2302 MUX2_X1 
XU1230 n563 n620 n500 n1208 NETTRAN_DUMMY_2303 NETTRAN_DUMMY_2304 MUX2_X1 
XU1229 n554 n543 n500 n1207 NETTRAN_DUMMY_2305 NETTRAN_DUMMY_2306 MUX2_X1 
XU1227 n1205 n1202 n453 n1206 NETTRAN_DUMMY_2307 NETTRAN_DUMMY_2308 MUX2_X1 
XU1226 n1204 n1203 n466 n1205 NETTRAN_DUMMY_2309 NETTRAN_DUMMY_2310 MUX2_X1 
XU1224 n620 n1763 n502 n1203 NETTRAN_DUMMY_2311 NETTRAN_DUMMY_2312 MUX2_X1 
XU1223 n1201 n1352 n502 n1202 NETTRAN_DUMMY_2313 NETTRAN_DUMMY_2314 MUX2_X1 
XU1222 n1791 n1752 n466 n1201 NETTRAN_DUMMY_2315 NETTRAN_DUMMY_2316 MUX2_X1 
XU1221 n1199 n1200 n433 d[30] NETTRAN_DUMMY_2317 NETTRAN_DUMMY_2318 MUX2_X1 
XU1219 n1198 n1193 n452 n1199 NETTRAN_DUMMY_2319 NETTRAN_DUMMY_2320 MUX2_X1 
XU1218 n1197 n1194 n445 n1198 NETTRAN_DUMMY_2321 NETTRAN_DUMMY_2322 MUX2_X1 
XU1217 n1196 n1195 n503 n1197 NETTRAN_DUMMY_2323 NETTRAN_DUMMY_2324 MUX2_X1 
XU1216 n615 n565 n473 n1196 NETTRAN_DUMMY_2325 NETTRAN_DUMMY_2326 MUX2_X1 
XU1215 n776 n1501 n473 n1195 NETTRAN_DUMMY_2327 NETTRAN_DUMMY_2328 MUX2_X1 
XU1214 n1671 n623 n503 n1194 NETTRAN_DUMMY_2329 NETTRAN_DUMMY_2330 MUX2_X1 
XU1213 n1191 n1192 n442 n1193 NETTRAN_DUMMY_2331 NETTRAN_DUMMY_2332 MUX2_X1 
XU1211 n1189 n1190 n503 n1191 NETTRAN_DUMMY_2333 NETTRAN_DUMMY_2334 MUX2_X1 
XU1209 n512 n1333 n473 n1189 NETTRAN_DUMMY_2335 NETTRAN_DUMMY_2336 MUX2_X1 
XU1208 n503 n1187 n445 n1188 NETTRAN_DUMMY_2337 NETTRAN_DUMMY_2338 MUX2_X1 
XU1206 n513 n1185 n452 n1186 NETTRAN_DUMMY_2339 NETTRAN_DUMMY_2340 MUX2_X1 
XU1205 n1184 n529 n445 n1185 NETTRAN_DUMMY_2341 NETTRAN_DUMMY_2342 MUX2_X1 
XU1204 n513 n569 n458 n1184 NETTRAN_DUMMY_2343 NETTRAN_DUMMY_2344 MUX2_X1 
XU1203 n1183 n1169 n433 d[2] NETTRAN_DUMMY_2345 NETTRAN_DUMMY_2346 MUX2_X1 
XU1202 n1182 n1176 n443 n1183 NETTRAN_DUMMY_2347 NETTRAN_DUMMY_2348 MUX2_X1 
XU1201 n1181 n1179 n455 n1182 NETTRAN_DUMMY_2349 NETTRAN_DUMMY_2350 MUX2_X1 
XU1200 n1180 n1806 n458 n1181 NETTRAN_DUMMY_2351 NETTRAN_DUMMY_2352 MUX2_X1 
XU1199 n606 n1499 n507 n1180 NETTRAN_DUMMY_2353 NETTRAN_DUMMY_2354 MUX2_X1 
XU1198 n1178 n1177 n458 n1179 NETTRAN_DUMMY_2355 NETTRAN_DUMMY_2356 MUX2_X1 
XU1197 n1742 n1749 n502 n1178 NETTRAN_DUMMY_2357 NETTRAN_DUMMY_2358 MUX2_X1 
XU1196 n493 n480 n495 n1177 NETTRAN_DUMMY_2359 NETTRAN_DUMMY_2360 MUX2_X1 
XU1195 n1175 n1172 n455 n1176 NETTRAN_DUMMY_2361 NETTRAN_DUMMY_2362 MUX2_X1 
XU1194 n1174 n1173 n471 n1175 NETTRAN_DUMMY_2363 NETTRAN_DUMMY_2364 MUX2_X1 
XU1193 n604 n583 n507 n1174 NETTRAN_DUMMY_2365 NETTRAN_DUMMY_2366 MUX2_X1 
XU1192 n1758 n1544 n502 n1173 NETTRAN_DUMMY_2367 NETTRAN_DUMMY_2368 MUX2_X1 
XU1191 n1170 n1171 n471 n1172 NETTRAN_DUMMY_2369 NETTRAN_DUMMY_2370 MUX2_X1 
XU1189 n549 n585 n502 n1170 NETTRAN_DUMMY_2371 NETTRAN_DUMMY_2372 MUX2_X1 
XU1188 n1168 n1161 n443 n1169 NETTRAN_DUMMY_2373 NETTRAN_DUMMY_2374 MUX2_X1 
XU1187 n1167 n1164 n455 n1168 NETTRAN_DUMMY_2375 NETTRAN_DUMMY_2376 MUX2_X1 
XU1186 n1165 n1166 n471 n1167 NETTRAN_DUMMY_2377 NETTRAN_DUMMY_2378 MUX2_X1 
XU1184 n1741 n582 n495 n1165 NETTRAN_DUMMY_2379 NETTRAN_DUMMY_2380 MUX2_X1 
XU1183 n1163 n1162 n471 n1164 NETTRAN_DUMMY_2381 NETTRAN_DUMMY_2382 MUX2_X1 
XU1182 n616 n551 n502 n1163 NETTRAN_DUMMY_2383 NETTRAN_DUMMY_2384 MUX2_X1 
XU1181 n587 n610 n502 n1162 NETTRAN_DUMMY_2385 NETTRAN_DUMMY_2386 MUX2_X1 
XU1180 n1158 n1159 n455 n1161 NETTRAN_DUMMY_2387 NETTRAN_DUMMY_2388 MUX2_X1 
XU1178 n1157 n1156 n471 n1158 NETTRAN_DUMMY_2389 NETTRAN_DUMMY_2390 MUX2_X1 
XU1177 n552 n1752 n502 n1157 NETTRAN_DUMMY_2391 NETTRAN_DUMMY_2392 MUX2_X1 
XU1176 n625 n1835 n502 n1156 NETTRAN_DUMMY_2393 NETTRAN_DUMMY_2394 MUX2_X1 
XU1175 n1155 n1141 n442 d[29] NETTRAN_DUMMY_2395 NETTRAN_DUMMY_2396 MUX2_X1 
XU1174 n1154 n1147 n452 n1155 NETTRAN_DUMMY_2397 NETTRAN_DUMMY_2398 MUX2_X1 
XU1173 n1153 n1150 n458 n1154 NETTRAN_DUMMY_2399 NETTRAN_DUMMY_2400 MUX2_X1 
XU1172 n1152 n1151 n495 n1153 NETTRAN_DUMMY_2401 NETTRAN_DUMMY_2402 MUX2_X1 
XU1171 n1812 n516 n433 n1152 NETTRAN_DUMMY_2403 NETTRAN_DUMMY_2404 MUX2_X1 
XU1170 n1530 n513 n433 n1151 NETTRAN_DUMMY_2405 NETTRAN_DUMMY_2406 MUX2_X1 
XU1169 n1149 n1148 n495 n1150 NETTRAN_DUMMY_2407 NETTRAN_DUMMY_2408 MUX2_X1 
XU1168 n594 n512 n433 n1149 NETTRAN_DUMMY_2409 NETTRAN_DUMMY_2410 MUX2_X1 
XU1167 n1819 n551 n435 n1148 NETTRAN_DUMMY_2411 NETTRAN_DUMMY_2412 MUX2_X1 
XU1166 n1146 n1144 n468 n1147 NETTRAN_DUMMY_2413 NETTRAN_DUMMY_2414 MUX2_X1 
XU1165 n1145 n546 n503 n1146 NETTRAN_DUMMY_2415 NETTRAN_DUMMY_2416 MUX2_X1 
XU1164 n1542 n512 n433 n1145 NETTRAN_DUMMY_2417 NETTRAN_DUMMY_2418 MUX2_X1 
XU1163 n1142 n1143 n503 n1144 NETTRAN_DUMMY_2419 NETTRAN_DUMMY_2420 MUX2_X1 
XU1161 n1832 n1500 n433 n1142 NETTRAN_DUMMY_2421 NETTRAN_DUMMY_2422 MUX2_X1 
XU1160 n1140 n1135 n452 n1141 NETTRAN_DUMMY_2423 NETTRAN_DUMMY_2424 MUX2_X1 
XU1159 n1139 n1138 n468 n1140 NETTRAN_DUMMY_2425 NETTRAN_DUMMY_2426 MUX2_X1 
XU1157 n1136 n1137 n503 n1138 NETTRAN_DUMMY_2427 NETTRAN_DUMMY_2428 MUX2_X1 
XU1155 n536 n1333 n433 n1136 NETTRAN_DUMMY_2429 NETTRAN_DUMMY_2430 MUX2_X1 
XU1154 n1134 n1132 n473 n1135 NETTRAN_DUMMY_2431 NETTRAN_DUMMY_2432 MUX2_X1 
XU1153 n513 n1133 n503 n1134 NETTRAN_DUMMY_2433 NETTRAN_DUMMY_2434 MUX2_X1 
XU1151 n1585 n431 n503 n1132 NETTRAN_DUMMY_2435 NETTRAN_DUMMY_2436 MUX2_X1 
XU1150 n1131 n1117 n435 d[28] NETTRAN_DUMMY_2437 NETTRAN_DUMMY_2438 MUX2_X1 
XU1149 n1130 n1123 n439 n1131 NETTRAN_DUMMY_2439 NETTRAN_DUMMY_2440 MUX2_X1 
XU1148 n1129 n1126 n452 n1130 NETTRAN_DUMMY_2441 NETTRAN_DUMMY_2442 MUX2_X1 
XU1147 n1128 n1127 n503 n1129 NETTRAN_DUMMY_2443 NETTRAN_DUMMY_2444 MUX2_X1 
XU1146 n516 n1768 n462 n1128 NETTRAN_DUMMY_2445 NETTRAN_DUMMY_2446 MUX2_X1 
XU1145 n533 n606 n462 n1127 NETTRAN_DUMMY_2447 NETTRAN_DUMMY_2448 MUX2_X1 
XU1144 n1125 n1124 n503 n1126 NETTRAN_DUMMY_2449 NETTRAN_DUMMY_2450 MUX2_X1 
XU1143 n590 n1789 n462 n1125 NETTRAN_DUMMY_2451 NETTRAN_DUMMY_2452 MUX2_X1 
XU1352 n1756 n488 n500 n1328 NETTRAN_DUMMY_2453 NETTRAN_DUMMY_2454 MUX2_X1 
XU1351 n1326 n1323 n453 n1327 NETTRAN_DUMMY_2455 NETTRAN_DUMMY_2456 MUX2_X1 
XU1350 n1325 n1324 n464 n1326 NETTRAN_DUMMY_2457 NETTRAN_DUMMY_2458 MUX2_X1 
XU1348 n626 n605 n500 n1324 NETTRAN_DUMMY_2459 NETTRAN_DUMMY_2460 MUX2_X1 
XU1347 n1321 n1322 n464 n1323 NETTRAN_DUMMY_2461 NETTRAN_DUMMY_2462 MUX2_X1 
XU1345 n595 n1748 n500 n1321 NETTRAN_DUMMY_2463 NETTRAN_DUMMY_2464 MUX2_X1 
XU1344 n1320 n1305 n435 d[38] NETTRAN_DUMMY_2465 NETTRAN_DUMMY_2466 MUX2_X1 
XU1343 n1319 n1312 n442 n1320 NETTRAN_DUMMY_2467 NETTRAN_DUMMY_2468 MUX2_X1 
XU1342 n13180 n1315 n453 n1319 NETTRAN_DUMMY_2469 NETTRAN_DUMMY_2470 MUX2_X1 
XU1341 n1317 n1316 n502 n13180 NETTRAN_DUMMY_2471 NETTRAN_DUMMY_2472 MUX2_X1 
XU1340 n578 n512 n466 n1317 NETTRAN_DUMMY_2473 NETTRAN_DUMMY_2474 MUX2_X1 
XU1339 n1842 n1799 n466 n1316 NETTRAN_DUMMY_2475 NETTRAN_DUMMY_2476 MUX2_X1 
XU1338 n1314 n1313 n502 n1315 NETTRAN_DUMMY_2477 NETTRAN_DUMMY_2478 MUX2_X1 
XU1337 n629 n612 n466 n1314 NETTRAN_DUMMY_2479 NETTRAN_DUMMY_2480 MUX2_X1 
XU1336 n1822 n584 n466 n1313 NETTRAN_DUMMY_2481 NETTRAN_DUMMY_2482 MUX2_X1 
XU1335 n1311 n1308 n453 n1312 NETTRAN_DUMMY_2483 NETTRAN_DUMMY_2484 MUX2_X1 
XU1334 n1309 n1310 n500 n1311 NETTRAN_DUMMY_2485 NETTRAN_DUMMY_2486 MUX2_X1 
XU1332 n558 n1522 n464 n1309 NETTRAN_DUMMY_2487 NETTRAN_DUMMY_2488 MUX2_X1 
XU1331 n1306 n1307 n500 n1308 NETTRAN_DUMMY_2489 NETTRAN_DUMMY_2490 MUX2_X1 
XU1329 n579 n578 n466 n1306 NETTRAN_DUMMY_2491 NETTRAN_DUMMY_2492 MUX2_X1 
XU1328 n1304 n1297 n442 n1305 NETTRAN_DUMMY_2493 NETTRAN_DUMMY_2494 MUX2_X1 
XU1327 n1303 n1301 n453 n1304 NETTRAN_DUMMY_2495 NETTRAN_DUMMY_2496 MUX2_X1 
XU1326 n1672 n1302 n500 n1303 NETTRAN_DUMMY_2497 NETTRAN_DUMMY_2498 MUX2_X1 
XU1325 n622 n593 n475 n1302 NETTRAN_DUMMY_2499 NETTRAN_DUMMY_2500 MUX2_X1 
XU1324 n1299 n1298 n500 n1301 NETTRAN_DUMMY_2501 NETTRAN_DUMMY_2502 MUX2_X1 
XU1322 n1523 n537 n475 n1298 NETTRAN_DUMMY_2503 NETTRAN_DUMMY_2504 MUX2_X1 
XU1321 n1296 n1292 n453 n1297 NETTRAN_DUMMY_2505 NETTRAN_DUMMY_2506 MUX2_X1 
XU1320 n1293 n1294 n500 n1296 NETTRAN_DUMMY_2507 NETTRAN_DUMMY_2508 MUX2_X1 
XU1318 n1766 n1816 n464 n1293 NETTRAN_DUMMY_2509 NETTRAN_DUMMY_2510 MUX2_X1 
XU1317 n1291 n1290 n500 n1292 NETTRAN_DUMMY_2511 NETTRAN_DUMMY_2512 MUX2_X1 
XU1315 n1545 n621 n464 n1290 NETTRAN_DUMMY_2513 NETTRAN_DUMMY_2514 MUX2_X1 
XU1314 n1289 n1274 n435 d[37] NETTRAN_DUMMY_2515 NETTRAN_DUMMY_2516 MUX2_X1 
XU1313 n1288 n1281 n442 n1289 NETTRAN_DUMMY_2517 NETTRAN_DUMMY_2518 MUX2_X1 
XU1312 n1287 n1284 n502 n1288 NETTRAN_DUMMY_2519 NETTRAN_DUMMY_2520 MUX2_X1 
XU1311 n1286 n1285 n466 n1287 NETTRAN_DUMMY_2521 NETTRAN_DUMMY_2522 MUX2_X1 
XU1309 n1751 n609 n453 n1285 NETTRAN_DUMMY_2523 NETTRAN_DUMMY_2524 MUX2_X1 
XU1308 n1283 n1282 n466 n1284 NETTRAN_DUMMY_2525 NETTRAN_DUMMY_2526 MUX2_X1 
XU1307 n579 n1754 n453 n1283 NETTRAN_DUMMY_2527 NETTRAN_DUMMY_2528 MUX2_X1 
XU1306 n1852 n1855 n453 n1282 NETTRAN_DUMMY_2529 NETTRAN_DUMMY_2530 MUX2_X1 
XU1305 n1280 n1277 n502 n1281 NETTRAN_DUMMY_2531 NETTRAN_DUMMY_2532 MUX2_X1 
XU1304 n1279 n1278 n466 n1280 NETTRAN_DUMMY_2533 NETTRAN_DUMMY_2534 MUX2_X1 
XU1303 n1842 n1832 n453 n1279 NETTRAN_DUMMY_2535 NETTRAN_DUMMY_2536 MUX2_X1 
XU1302 n493 n552 n453 n1278 NETTRAN_DUMMY_2537 NETTRAN_DUMMY_2538 MUX2_X1 
XU1301 n1276 n1275 n466 n1277 NETTRAN_DUMMY_2539 NETTRAN_DUMMY_2540 MUX2_X1 
XU1299 n612 n1758 n453 n1275 NETTRAN_DUMMY_2541 NETTRAN_DUMMY_2542 MUX2_X1 
XU1298 n1273 n1266 n442 n1274 NETTRAN_DUMMY_2543 NETTRAN_DUMMY_2544 MUX2_X1 
XU1297 n1272 n1269 n500 n1273 NETTRAN_DUMMY_2545 NETTRAN_DUMMY_2546 MUX2_X1 
XU1296 n1271 n1270 n464 n1272 NETTRAN_DUMMY_2547 NETTRAN_DUMMY_2548 MUX2_X1 
XU1295 n1530 n560 n453 n1271 NETTRAN_DUMMY_2549 NETTRAN_DUMMY_2550 MUX2_X1 
XU1294 n1523 n1828 n453 n1270 NETTRAN_DUMMY_2551 NETTRAN_DUMMY_2552 MUX2_X1 
XU1293 n1268 n1267 n466 n1269 NETTRAN_DUMMY_2553 NETTRAN_DUMMY_2554 MUX2_X1 
XU1292 n1742 n520 n453 n1268 NETTRAN_DUMMY_2555 NETTRAN_DUMMY_2556 MUX2_X1 
XU1291 n1767 n1805 n453 n1267 NETTRAN_DUMMY_2557 NETTRAN_DUMMY_2558 MUX2_X1 
XU1290 n1265 n1262 n500 n1266 NETTRAN_DUMMY_2559 NETTRAN_DUMMY_2560 MUX2_X1 
XU1289 n1264 n1263 n466 n1265 NETTRAN_DUMMY_2561 NETTRAN_DUMMY_2562 MUX2_X1 
XU1288 n1756 n1772 n453 n1264 NETTRAN_DUMMY_2563 NETTRAN_DUMMY_2564 MUX2_X1 
XU1287 n554 n1543 n453 n1263 NETTRAN_DUMMY_2565 NETTRAN_DUMMY_2566 MUX2_X1 
XU1286 n1261 n1260 n466 n1262 NETTRAN_DUMMY_2567 NETTRAN_DUMMY_2568 MUX2_X1 
XU1285 n1827 n625 n453 n1261 NETTRAN_DUMMY_2569 NETTRAN_DUMMY_2570 MUX2_X1 
XU1284 n1841 n1752 n453 n1260 NETTRAN_DUMMY_2571 NETTRAN_DUMMY_2572 MUX2_X1 
XU1283 n1259 n1243 n435 d[36] NETTRAN_DUMMY_2573 NETTRAN_DUMMY_2574 MUX2_X1 
XU1282 n1258 n1250 n443 n1259 NETTRAN_DUMMY_2575 NETTRAN_DUMMY_2576 MUX2_X1 
XU1281 n1257 n1253 n453 n1258 NETTRAN_DUMMY_2577 NETTRAN_DUMMY_2578 MUX2_X1 
XU1280 n1256 n1254 n466 n1257 NETTRAN_DUMMY_2579 NETTRAN_DUMMY_2580 MUX2_X1 
XU1279 n526 n1255 n509 n1256 NETTRAN_DUMMY_2581 NETTRAN_DUMMY_2582 MUX2_X1 
XU1278 n528 n480 n495 n1255 NETTRAN_DUMMY_2583 NETTRAN_DUMMY_2584 MUX2_X1 
XU1277 n1835 n559 n502 n1254 NETTRAN_DUMMY_2585 NETTRAN_DUMMY_2586 MUX2_X1 
XU1276 n1252 n1251 n466 n1253 NETTRAN_DUMMY_2587 NETTRAN_DUMMY_2588 MUX2_X1 
XU1275 n1852 n611 n502 n1252 NETTRAN_DUMMY_2589 NETTRAN_DUMMY_2590 MUX2_X1 
XU1274 n612 n1753 n502 n1251 NETTRAN_DUMMY_2591 NETTRAN_DUMMY_2592 MUX2_X1 
XU1273 n1249 n1246 n453 n1250 NETTRAN_DUMMY_2593 NETTRAN_DUMMY_2594 MUX2_X1 
XU1272 n1248 n1247 n466 n1249 NETTRAN_DUMMY_2595 NETTRAN_DUMMY_2596 MUX2_X1 
XU1271 n1805 n603 n502 n1248 NETTRAN_DUMMY_2597 NETTRAN_DUMMY_2598 MUX2_X1 
XU1270 n1770 n607 n502 n1247 NETTRAN_DUMMY_2599 NETTRAN_DUMMY_2600 MUX2_X1 
XU1269 n1245 n1244 n466 n1246 NETTRAN_DUMMY_2601 NETTRAN_DUMMY_2602 MUX2_X1 
XU1268 n1747 n1774 n502 n1245 NETTRAN_DUMMY_2603 NETTRAN_DUMMY_2604 MUX2_X1 
XU1267 n541 n577 n502 n1244 NETTRAN_DUMMY_2605 NETTRAN_DUMMY_2606 MUX2_X1 
XU1266 n1242 n1235 n443 n1243 NETTRAN_DUMMY_2607 NETTRAN_DUMMY_2608 MUX2_X1 
XU1265 n1241 n1238 n453 n1242 NETTRAN_DUMMY_2609 NETTRAN_DUMMY_2610 MUX2_X1 
XU1264 n1240 n1239 n466 n1241 NETTRAN_DUMMY_2611 NETTRAN_DUMMY_2612 MUX2_X1 
XU1263 n532 n589 n502 n1240 NETTRAN_DUMMY_2613 NETTRAN_DUMMY_2614 MUX2_X1 
XU1262 n609 n536 n502 n1239 NETTRAN_DUMMY_2615 NETTRAN_DUMMY_2616 MUX2_X1 
XU1261 n1237 n1236 n466 n1238 NETTRAN_DUMMY_2617 NETTRAN_DUMMY_2618 MUX2_X1 
XU1260 n1752 n1797 n502 n1237 NETTRAN_DUMMY_2619 NETTRAN_DUMMY_2620 MUX2_X1 
XU1259 n1814 n1775 n502 n1236 NETTRAN_DUMMY_2621 NETTRAN_DUMMY_2622 MUX2_X1 
XU1258 n1234 n1231 n453 n1235 NETTRAN_DUMMY_2623 NETTRAN_DUMMY_2624 MUX2_X1 
XU1257 n1233 n1232 n466 n1234 NETTRAN_DUMMY_2625 NETTRAN_DUMMY_2626 MUX2_X1 
XU1256 n1824 n1544 n502 n1233 NETTRAN_DUMMY_2627 NETTRAN_DUMMY_2628 MUX2_X1 
XU1255 n1826 n610 n502 n1232 NETTRAN_DUMMY_2629 NETTRAN_DUMMY_2630 MUX2_X1 
XU1254 n1230 n1229 n466 n1231 NETTRAN_DUMMY_2631 NETTRAN_DUMMY_2632 MUX2_X1 
XU1251 n1228 n1214 n435 d[35] NETTRAN_DUMMY_2633 NETTRAN_DUMMY_2634 MUX2_X1 
XU1250 n1227 n1221 n442 n1228 NETTRAN_DUMMY_2635 NETTRAN_DUMMY_2636 MUX2_X1 
XU1249 n1226 n1224 n453 n1227 NETTRAN_DUMMY_2637 NETTRAN_DUMMY_2638 MUX2_X1 
XU1451 n595 n515 n477 n1426 NETTRAN_DUMMY_2639 NETTRAN_DUMMY_2640 MUX2_X1 
XU1450 n1761 n601 n477 n1425 NETTRAN_DUMMY_2641 NETTRAN_DUMMY_2642 MUX2_X1 
XU1449 n1423 n1416 n439 n1424 NETTRAN_DUMMY_2643 NETTRAN_DUMMY_2644 MUX2_X1 
XU1448 n1422 n1419 n454 n1423 NETTRAN_DUMMY_2645 NETTRAN_DUMMY_2646 MUX2_X1 
XU1447 n1421 n1420 n500 n1422 NETTRAN_DUMMY_2647 NETTRAN_DUMMY_2648 MUX2_X1 
XU1446 n1752 n621 n464 n1421 NETTRAN_DUMMY_2649 NETTRAN_DUMMY_2650 MUX2_X1 
XU1445 n517 n1850 n464 n1420 NETTRAN_DUMMY_2651 NETTRAN_DUMMY_2652 MUX2_X1 
XU1444 n1418 n1417 n499 n1419 NETTRAN_DUMMY_2653 NETTRAN_DUMMY_2654 MUX2_X1 
XU1443 n1832 n1761 n477 n1418 NETTRAN_DUMMY_2655 NETTRAN_DUMMY_2656 MUX2_X1 
XU1442 n515 n590 n477 n1417 NETTRAN_DUMMY_2657 NETTRAN_DUMMY_2658 MUX2_X1 
XU1441 n1415 n1412 n454 n1416 NETTRAN_DUMMY_2659 NETTRAN_DUMMY_2660 MUX2_X1 
XU1440 n1414 n1413 n499 n1415 NETTRAN_DUMMY_2661 NETTRAN_DUMMY_2662 MUX2_X1 
XU1439 n1529 n564 n477 n1414 NETTRAN_DUMMY_2663 NETTRAN_DUMMY_2664 MUX2_X1 
XU1438 n516 n1530 n477 n1413 NETTRAN_DUMMY_2665 NETTRAN_DUMMY_2666 MUX2_X1 
XU1437 n1411 n1410 n499 n1412 NETTRAN_DUMMY_2667 NETTRAN_DUMMY_2668 MUX2_X1 
XU1435 n536 n621 n464 n1410 NETTRAN_DUMMY_2669 NETTRAN_DUMMY_2670 MUX2_X1 
XU1434 n1409 n1395 n435 d[40] NETTRAN_DUMMY_2671 NETTRAN_DUMMY_2672 MUX2_X1 
XU1433 n1408 n1402 n442 n1409 NETTRAN_DUMMY_2673 NETTRAN_DUMMY_2674 MUX2_X1 
XU1432 n1407 n1404 n454 n1408 NETTRAN_DUMMY_2675 NETTRAN_DUMMY_2676 MUX2_X1 
XU1431 n1406 n1405 n477 n1407 NETTRAN_DUMMY_2677 NETTRAN_DUMMY_2678 MUX2_X1 
XU1429 n526 n601 n499 n1405 NETTRAN_DUMMY_2679 NETTRAN_DUMMY_2680 MUX2_X1 
XU1428 n1850 n1403 n428 n1404 NETTRAN_DUMMY_2681 NETTRAN_DUMMY_2682 MUX2_X1 
XU1427 n1797 n1801 n471 n1403 NETTRAN_DUMMY_2683 NETTRAN_DUMMY_2684 MUX2_X1 
XU1426 n1401 n1398 n454 n1402 NETTRAN_DUMMY_2685 NETTRAN_DUMMY_2686 MUX2_X1 
XU1425 n1400 n1399 n477 n1401 NETTRAN_DUMMY_2687 NETTRAN_DUMMY_2688 MUX2_X1 
XU1424 n608 n1352 n499 n1400 NETTRAN_DUMMY_2689 NETTRAN_DUMMY_2690 MUX2_X1 
XU1423 n564 n596 n499 n1399 NETTRAN_DUMMY_2691 NETTRAN_DUMMY_2692 MUX2_X1 
XU1422 n1397 n1396 n477 n1398 NETTRAN_DUMMY_2693 NETTRAN_DUMMY_2694 MUX2_X1 
XU1421 n611 n581 n499 n1397 NETTRAN_DUMMY_2695 NETTRAN_DUMMY_2696 MUX2_X1 
XU1420 n526 n1765 n500 n1396 NETTRAN_DUMMY_2697 NETTRAN_DUMMY_2698 MUX2_X1 
XU1419 n1394 n1387 n442 n1395 NETTRAN_DUMMY_2699 NETTRAN_DUMMY_2700 MUX2_X1 
XU1418 n1393 n1390 n453 n1394 NETTRAN_DUMMY_2701 NETTRAN_DUMMY_2702 MUX2_X1 
XU1417 n1392 n1391 n464 n1393 NETTRAN_DUMMY_2703 NETTRAN_DUMMY_2704 MUX2_X1 
XU1416 n586 n599 n500 n1392 NETTRAN_DUMMY_2705 NETTRAN_DUMMY_2706 MUX2_X1 
XU1415 n548 n1774 n500 n1391 NETTRAN_DUMMY_2707 NETTRAN_DUMMY_2708 MUX2_X1 
XU1414 n1389 n1388 n464 n1390 NETTRAN_DUMMY_2709 NETTRAN_DUMMY_2710 MUX2_X1 
XU1413 n543 n1756 n500 n1389 NETTRAN_DUMMY_2711 NETTRAN_DUMMY_2712 MUX2_X1 
XU1412 n1771 n1318 n500 n1388 NETTRAN_DUMMY_2713 NETTRAN_DUMMY_2714 MUX2_X1 
XU1411 n1386 n1383 n453 n1387 NETTRAN_DUMMY_2715 NETTRAN_DUMMY_2716 MUX2_X1 
XU1410 n1385 n1384 n464 n1386 NETTRAN_DUMMY_2717 NETTRAN_DUMMY_2718 MUX2_X1 
XU1409 n528 n520 n500 n1385 NETTRAN_DUMMY_2719 NETTRAN_DUMMY_2720 MUX2_X1 
XU1408 n578 n616 n500 n1384 NETTRAN_DUMMY_2721 NETTRAN_DUMMY_2722 MUX2_X1 
XU1407 n1382 n1381 n464 n1383 NETTRAN_DUMMY_2723 NETTRAN_DUMMY_2724 MUX2_X1 
XU1406 n543 n1541 n500 n1382 NETTRAN_DUMMY_2725 NETTRAN_DUMMY_2726 MUX2_X1 
XU1405 n618 n1352 n500 n1381 NETTRAN_DUMMY_2727 NETTRAN_DUMMY_2728 MUX2_X1 
XU1404 n1380 n1363 n433 d[3] NETTRAN_DUMMY_2729 NETTRAN_DUMMY_2730 MUX2_X1 
XU1403 n1379 n1372 n443 n1380 NETTRAN_DUMMY_2731 NETTRAN_DUMMY_2732 MUX2_X1 
XU1402 n1378 n1375 n453 n1379 NETTRAN_DUMMY_2733 NETTRAN_DUMMY_2734 MUX2_X1 
XU1401 n1377 n1376 n471 n1378 NETTRAN_DUMMY_2735 NETTRAN_DUMMY_2736 MUX2_X1 
XU1400 n523 n620 n502 n1377 NETTRAN_DUMMY_2737 NETTRAN_DUMMY_2738 MUX2_X1 
XU1399 n562 n1776 n502 n1376 NETTRAN_DUMMY_2739 NETTRAN_DUMMY_2740 MUX2_X1 
XU1398 n1374 n1373 n471 n1375 NETTRAN_DUMMY_2741 NETTRAN_DUMMY_2742 MUX2_X1 
XU1397 n1539 n1751 n502 n1374 NETTRAN_DUMMY_2743 NETTRAN_DUMMY_2744 MUX2_X1 
XU1396 n569 n561 n502 n1373 NETTRAN_DUMMY_2745 NETTRAN_DUMMY_2746 MUX2_X1 
XU1395 n1371 n1367 n453 n1372 NETTRAN_DUMMY_2747 NETTRAN_DUMMY_2748 MUX2_X1 
XU1394 n1370 n1368 n475 n1371 NETTRAN_DUMMY_2749 NETTRAN_DUMMY_2750 MUX2_X1 
XU1393 n593 n1369 n502 n1370 NETTRAN_DUMMY_2751 NETTRAN_DUMMY_2752 MUX2_X1 
XU1391 n1746 n605 n507 n1368 NETTRAN_DUMMY_2753 NETTRAN_DUMMY_2754 MUX2_X1 
XU1390 n1365 n1364 n471 n1367 NETTRAN_DUMMY_2755 NETTRAN_DUMMY_2756 MUX2_X1 
XU1388 n1805 n1808 n502 n1364 NETTRAN_DUMMY_2757 NETTRAN_DUMMY_2758 MUX2_X1 
XU1387 n1362 n1355 n443 n1363 NETTRAN_DUMMY_2759 NETTRAN_DUMMY_2760 MUX2_X1 
XU1386 n1361 n1358 n453 n1362 NETTRAN_DUMMY_2761 NETTRAN_DUMMY_2762 MUX2_X1 
XU1385 n1360 n1359 n466 n1361 NETTRAN_DUMMY_2763 NETTRAN_DUMMY_2764 MUX2_X1 
XU1384 n1814 n550 n502 n1360 NETTRAN_DUMMY_2765 NETTRAN_DUMMY_2766 MUX2_X1 
XU1383 n1500 n620 n502 n1359 NETTRAN_DUMMY_2767 NETTRAN_DUMMY_2768 MUX2_X1 
XU1382 n1357 n1356 n475 n1358 NETTRAN_DUMMY_2769 NETTRAN_DUMMY_2770 MUX2_X1 
XU1381 n1352 n1674 n507 n1357 NETTRAN_DUMMY_2771 NETTRAN_DUMMY_2772 MUX2_X1 
XU1380 n547 n1746 n507 n1356 NETTRAN_DUMMY_2773 NETTRAN_DUMMY_2774 MUX2_X1 
XU1379 n13520 n1353 n453 n1355 NETTRAN_DUMMY_2775 NETTRAN_DUMMY_2776 MUX2_X1 
XU1377 n1351 n1350 n466 n13520 NETTRAN_DUMMY_2777 NETTRAN_DUMMY_2778 MUX2_X1 
XU1376 n1754 n1745 n502 n1351 NETTRAN_DUMMY_2779 NETTRAN_DUMMY_2780 MUX2_X1 
XU1375 n611 n1776 n502 n1350 NETTRAN_DUMMY_2781 NETTRAN_DUMMY_2782 MUX2_X1 
XU1374 n1349 n1335 n435 d[39] NETTRAN_DUMMY_2783 NETTRAN_DUMMY_2784 MUX2_X1 
XU1373 n1348 n1342 n442 n1349 NETTRAN_DUMMY_2785 NETTRAN_DUMMY_2786 MUX2_X1 
XU1372 n1347 n1344 n453 n1348 NETTRAN_DUMMY_2787 NETTRAN_DUMMY_2788 MUX2_X1 
XU1371 n1346 n1345 n466 n1347 NETTRAN_DUMMY_2789 NETTRAN_DUMMY_2790 MUX2_X1 
XU1370 n598 n540 n500 n1346 NETTRAN_DUMMY_2791 NETTRAN_DUMMY_2792 MUX2_X1 
XU1369 n1827 n1745 n502 n1345 NETTRAN_DUMMY_2793 NETTRAN_DUMMY_2794 MUX2_X1 
XU1368 n1757 n1343 n466 n1344 NETTRAN_DUMMY_2795 NETTRAN_DUMMY_2796 MUX2_X1 
XU1367 n1845 n1826 n500 n1343 NETTRAN_DUMMY_2797 NETTRAN_DUMMY_2798 MUX2_X1 
XU1366 n1341 n1338 n453 n1342 NETTRAN_DUMMY_2799 NETTRAN_DUMMY_2800 MUX2_X1 
XU1365 n1340 n1339 n466 n1341 NETTRAN_DUMMY_2801 NETTRAN_DUMMY_2802 MUX2_X1 
XU1364 n552 n618 n502 n1340 NETTRAN_DUMMY_2803 NETTRAN_DUMMY_2804 MUX2_X1 
XU1363 n527 n1535 n507 n1339 NETTRAN_DUMMY_2805 NETTRAN_DUMMY_2806 MUX2_X1 
XU1362 n1337 n1336 n466 n1338 NETTRAN_DUMMY_2807 NETTRAN_DUMMY_2808 MUX2_X1 
XU1360 n1544 n1796 n502 n1336 NETTRAN_DUMMY_2809 NETTRAN_DUMMY_2810 MUX2_X1 
XU1359 n1334 n1327 n442 n1335 NETTRAN_DUMMY_2811 NETTRAN_DUMMY_2812 MUX2_X1 
XU1358 n13330 n1330 n453 n1334 NETTRAN_DUMMY_2813 NETTRAN_DUMMY_2814 MUX2_X1 
XU1357 n1332 n1331 n464 n13330 NETTRAN_DUMMY_2815 NETTRAN_DUMMY_2816 MUX2_X1 
XU1356 n625 n529 n500 n1332 NETTRAN_DUMMY_2817 NETTRAN_DUMMY_2818 MUX2_X1 
XU1355 n570 n1318 n500 n1331 NETTRAN_DUMMY_2819 NETTRAN_DUMMY_2820 MUX2_X1 
XU1354 n1329 n1328 n464 n1330 NETTRAN_DUMMY_2821 NETTRAN_DUMMY_2822 MUX2_X1 
XU1353 n1819 n1841 n500 n1329 NETTRAN_DUMMY_2823 NETTRAN_DUMMY_2824 MUX2_X1 
XU1557 n1520 n488 n509 n1515 NETTRAN_DUMMY_2825 NETTRAN_DUMMY_2826 MUX2_X1 
XU1556 n1513 n1514 n452 n1116 NETTRAN_DUMMY_2827 NETTRAN_DUMMY_2828 MUX2_X1 
XU1554 n512 n593 n473 n1513 NETTRAN_DUMMY_2829 NETTRAN_DUMMY_2830 MUX2_X1 
XU1553 n1525 n1318 n509 n1512 NETTRAN_DUMMY_2831 NETTRAN_DUMMY_2832 MUX2_X1 
XU1552 n628 n1528 n499 n1084 NETTRAN_DUMMY_2833 NETTRAN_DUMMY_2834 MUX2_X1 
XU1551 n492 n1760 n475 n1511 NETTRAN_DUMMY_2835 NETTRAN_DUMMY_2836 MUX2_X1 
XU1550 n560 n1538 n507 n1027 NETTRAN_DUMMY_2837 NETTRAN_DUMMY_2838 MUX2_X1 
XU1549 n526 n517 n509 n1510 NETTRAN_DUMMY_2839 NETTRAN_DUMMY_2840 MUX2_X1 
XU1548 n493 n1526 n509 n1509 NETTRAN_DUMMY_2841 NETTRAN_DUMMY_2842 MUX2_X1 
XU1547 n604 n1535 n507 n1508 NETTRAN_DUMMY_2843 NETTRAN_DUMMY_2844 MUX2_X1 
XU1546 n492 n488 n515 n1507 NETTRAN_DUMMY_2845 NETTRAN_DUMMY_2846 MUX2_X1 
XU1545 n1333 n628 n497 n884 NETTRAN_DUMMY_2847 NETTRAN_DUMMY_2848 MUX2_X1 
XU1544 n1840 n572 n507 n855 NETTRAN_DUMMY_2849 NETTRAN_DUMMY_2850 MUX2_X1 
XU1543 n526 n493 n509 n1506 NETTRAN_DUMMY_2851 NETTRAN_DUMMY_2852 MUX2_X1 
XU1542 n488 n1520 n509 n1505 NETTRAN_DUMMY_2853 NETTRAN_DUMMY_2854 MUX2_X1 
XU1541 n1522 n1816 n507 n765 NETTRAN_DUMMY_2855 NETTRAN_DUMMY_2856 MUX2_X1 
XU1540 n516 n1543 n473 n1504 NETTRAN_DUMMY_2857 NETTRAN_DUMMY_2858 MUX2_X1 
XU1539 n513 n525 n468 n734 NETTRAN_DUMMY_2859 NETTRAN_DUMMY_2860 MUX2_X1 
XU1538 n627 n1501 n473 n1503 NETTRAN_DUMMY_2861 NETTRAN_DUMMY_2862 MUX2_X1 
XU1537 n513 n1498 n448 n1502 NETTRAN_DUMMY_2863 NETTRAN_DUMMY_2864 MUX2_X1 
XU1526 n528 n488 n515 n1497 NETTRAN_DUMMY_2865 NETTRAN_DUMMY_2866 MUX2_X1 
XU1525 n615 n462 n1070 NETTRAN_DUMMY_2867 NETTRAN_DUMMY_2868 XOR2_X1 
XU1524 n1496 n1482 n435 d[43] NETTRAN_DUMMY_2869 NETTRAN_DUMMY_2870 MUX2_X1 
XU1523 n1495 n1488 n439 n1496 NETTRAN_DUMMY_2871 NETTRAN_DUMMY_2872 MUX2_X1 
XU1522 n1494 n1491 n454 n1495 NETTRAN_DUMMY_2873 NETTRAN_DUMMY_2874 MUX2_X1 
XU1521 n1493 n1492 n499 n1494 NETTRAN_DUMMY_2875 NETTRAN_DUMMY_2876 MUX2_X1 
XU1520 n1811 n605 n477 n1493 NETTRAN_DUMMY_2877 NETTRAN_DUMMY_2878 MUX2_X1 
XU1519 n553 n577 n477 n1492 NETTRAN_DUMMY_2879 NETTRAN_DUMMY_2880 MUX2_X1 
XU1518 n1490 n1489 n499 n1491 NETTRAN_DUMMY_2881 NETTRAN_DUMMY_2882 MUX2_X1 
XU1517 n563 n1541 n477 n1490 NETTRAN_DUMMY_2883 NETTRAN_DUMMY_2884 MUX2_X1 
XU1516 n1761 n1533 n477 n1489 NETTRAN_DUMMY_2885 NETTRAN_DUMMY_2886 MUX2_X1 
XU1515 n1487 n1485 n454 n1488 NETTRAN_DUMMY_2887 NETTRAN_DUMMY_2888 MUX2_X1 
XU1514 n1673 n1486 n499 n1487 NETTRAN_DUMMY_2889 NETTRAN_DUMMY_2890 MUX2_X1 
XU1513 n1520 n488 n477 n1486 NETTRAN_DUMMY_2891 NETTRAN_DUMMY_2892 MUX2_X1 
XU1512 n1484 n1483 n499 n1485 NETTRAN_DUMMY_2893 NETTRAN_DUMMY_2894 MUX2_X1 
XU1511 n1787 n492 n477 n1484 NETTRAN_DUMMY_2895 NETTRAN_DUMMY_2896 MUX2_X1 
XU1510 n1542 n564 n477 n1483 NETTRAN_DUMMY_2897 NETTRAN_DUMMY_2898 MUX2_X1 
XU1509 n1481 n1474 n439 n1482 NETTRAN_DUMMY_2899 NETTRAN_DUMMY_2900 MUX2_X1 
XU1508 n1480 n1477 n454 n1481 NETTRAN_DUMMY_2901 NETTRAN_DUMMY_2902 MUX2_X1 
XU1507 n1479 n1478 n499 n1480 NETTRAN_DUMMY_2903 NETTRAN_DUMMY_2904 MUX2_X1 
XU1506 n1773 IN1 n462 n1479 NETTRAN_DUMMY_2905 NETTRAN_DUMMY_2906 MUX2_X1 
XU1505 n1755 n612 n462 n1478 NETTRAN_DUMMY_2907 NETTRAN_DUMMY_2908 MUX2_X1 
XU1504 n1476 n1475 n499 n1477 NETTRAN_DUMMY_2909 NETTRAN_DUMMY_2910 MUX2_X1 
XU1503 n535 n1318 n462 n1476 NETTRAN_DUMMY_2911 NETTRAN_DUMMY_2912 MUX2_X1 
XU1502 n516 n567 n462 n1475 NETTRAN_DUMMY_2913 NETTRAN_DUMMY_2914 MUX2_X1 
XU1501 n1473 n1470 n454 n1474 NETTRAN_DUMMY_2915 NETTRAN_DUMMY_2916 MUX2_X1 
XU1500 n1472 n1471 n499 n1473 NETTRAN_DUMMY_2917 NETTRAN_DUMMY_2918 MUX2_X1 
XU1499 n533 n1523 n477 n1472 NETTRAN_DUMMY_2919 NETTRAN_DUMMY_2920 MUX2_X1 
XU1498 n579 n1533 n477 n1471 NETTRAN_DUMMY_2921 NETTRAN_DUMMY_2922 MUX2_X1 
XU1497 n1469 n1673 n499 n1470 NETTRAN_DUMMY_2923 NETTRAN_DUMMY_2924 MUX2_X1 
XU1496 n493 n488 n477 n1469 NETTRAN_DUMMY_2925 NETTRAN_DUMMY_2926 MUX2_X1 
XU1495 n1468 n1454 n435 d[42] NETTRAN_DUMMY_2927 NETTRAN_DUMMY_2928 MUX2_X1 
XU1494 n1467 n1460 n442 n1468 NETTRAN_DUMMY_2929 NETTRAN_DUMMY_2930 MUX2_X1 
XU1493 n1466 n1463 n453 n1467 NETTRAN_DUMMY_2931 NETTRAN_DUMMY_2932 MUX2_X1 
XU1492 n1465 n1464 n500 n1466 NETTRAN_DUMMY_2933 NETTRAN_DUMMY_2934 MUX2_X1 
XU1491 n545 n1847 n464 n1465 NETTRAN_DUMMY_2935 NETTRAN_DUMMY_2936 MUX2_X1 
XU1490 n523 n1852 n464 n1464 NETTRAN_DUMMY_2937 NETTRAN_DUMMY_2938 MUX2_X1 
XU1489 n1462 n1461 n500 n1463 NETTRAN_DUMMY_2939 NETTRAN_DUMMY_2940 MUX2_X1 
XU1488 n1832 n593 n464 n1462 NETTRAN_DUMMY_2941 NETTRAN_DUMMY_2942 MUX2_X1 
XU1487 n1525 n540 n464 n1461 NETTRAN_DUMMY_2943 NETTRAN_DUMMY_2944 MUX2_X1 
XU1486 n1459 n1457 n453 n1460 NETTRAN_DUMMY_2945 NETTRAN_DUMMY_2946 MUX2_X1 
XU1485 n1458 n633 n500 n1459 NETTRAN_DUMMY_2947 NETTRAN_DUMMY_2948 MUX2_X1 
XU1484 n526 n612 n464 n1458 NETTRAN_DUMMY_2949 NETTRAN_DUMMY_2950 MUX2_X1 
XU1483 n1456 n1455 n500 n1457 NETTRAN_DUMMY_2951 NETTRAN_DUMMY_2952 MUX2_X1 
XU1482 n1797 n516 n466 n1456 NETTRAN_DUMMY_2953 NETTRAN_DUMMY_2954 MUX2_X1 
XU1481 n1773 n612 n464 n1455 NETTRAN_DUMMY_2955 NETTRAN_DUMMY_2956 MUX2_X1 
XU1480 n1453 n1446 n442 n1454 NETTRAN_DUMMY_2957 NETTRAN_DUMMY_2958 MUX2_X1 
XU1479 n1452 n1449 n454 n1453 NETTRAN_DUMMY_2959 NETTRAN_DUMMY_2960 MUX2_X1 
XU1478 n1451 n1450 n500 n1452 NETTRAN_DUMMY_2961 NETTRAN_DUMMY_2962 MUX2_X1 
XU1477 n530 n618 n464 n1451 NETTRAN_DUMMY_2963 NETTRAN_DUMMY_2964 MUX2_X1 
XU1476 n1844 n1533 n464 n1450 NETTRAN_DUMMY_2965 NETTRAN_DUMMY_2966 MUX2_X1 
XU1475 n1448 n1447 n500 n1449 NETTRAN_DUMMY_2967 NETTRAN_DUMMY_2968 MUX2_X1 
XU1473 n516 n530 n477 n1447 NETTRAN_DUMMY_2969 NETTRAN_DUMMY_2970 MUX2_X1 
XU1472 n1445 n1442 n454 n1446 NETTRAN_DUMMY_2971 NETTRAN_DUMMY_2972 MUX2_X1 
XU1471 n1444 n1443 n500 n1445 NETTRAN_DUMMY_2973 NETTRAN_DUMMY_2974 MUX2_X1 
XU1470 n584 n1833 n464 n1444 NETTRAN_DUMMY_2975 NETTRAN_DUMMY_2976 MUX2_X1 
XU1469 n493 n554 n464 n1443 NETTRAN_DUMMY_2977 NETTRAN_DUMMY_2978 MUX2_X1 
XU1468 n1441 n1440 n500 n1442 NETTRAN_DUMMY_2979 NETTRAN_DUMMY_2980 MUX2_X1 
XU1467 n515 n585 n464 n1441 NETTRAN_DUMMY_2981 NETTRAN_DUMMY_2982 MUX2_X1 
XU1466 n1538 n1543 n464 n1440 NETTRAN_DUMMY_2983 NETTRAN_DUMMY_2984 MUX2_X1 
XU1465 n1439 n1424 n435 d[41] NETTRAN_DUMMY_2985 NETTRAN_DUMMY_2986 MUX2_X1 
XU1464 n1438 n1431 n439 n1439 NETTRAN_DUMMY_2987 NETTRAN_DUMMY_2988 MUX2_X1 
XU1463 n1437 n1434 n454 n1438 NETTRAN_DUMMY_2989 NETTRAN_DUMMY_2990 MUX2_X1 
XU1462 n1436 n1435 n499 n1437 NETTRAN_DUMMY_2991 NETTRAN_DUMMY_2992 MUX2_X1 
XU1461 n1545 n605 n477 n1436 NETTRAN_DUMMY_2993 NETTRAN_DUMMY_2994 MUX2_X1 
XU1460 n531 n1815 n477 n1435 NETTRAN_DUMMY_2995 NETTRAN_DUMMY_2996 MUX2_X1 
XU1459 n1433 n1432 n499 n1434 NETTRAN_DUMMY_2997 NETTRAN_DUMMY_2998 MUX2_X1 
XU1458 n1529 n1766 n477 n1433 NETTRAN_DUMMY_2999 NETTRAN_DUMMY_3000 MUX2_X1 
XU1457 n760 n611 n477 n1432 NETTRAN_DUMMY_3001 NETTRAN_DUMMY_3002 MUX2_X1 
XU1456 n1430 n1427 n454 n1431 NETTRAN_DUMMY_3003 NETTRAN_DUMMY_3004 MUX2_X1 
XU1455 n1428 n1429 n499 n1430 NETTRAN_DUMMY_3005 NETTRAN_DUMMY_3006 MUX2_X1 
XU1453 n535 n575 n477 n1428 NETTRAN_DUMMY_3007 NETTRAN_DUMMY_3008 MUX2_X1 
XU1452 n1426 n1425 n499 n1427 NETTRAN_DUMMY_3009 NETTRAN_DUMMY_3010 MUX2_X1 
XU450 n622 n1827 NETTRAN_DUMMY_3011 NETTRAN_DUMMY_3012 INV_X1 
XU449 n556 n1835 NETTRAN_DUMMY_3013 NETTRAN_DUMMY_3014 INV_X1 
XU448 n21 n1617 NETTRAN_DUMMY_3015 NETTRAN_DUMMY_3016 INV_X1 
XU447 n545 n1766 NETTRAN_DUMMY_3017 NETTRAN_DUMMY_3018 INV_X1 
XU446 n750 n1669 NETTRAN_DUMMY_3019 NETTRAN_DUMMY_3020 INV_X1 
XU445 n43 n1634 NETTRAN_DUMMY_3021 NETTRAN_DUMMY_3022 INV_X1 
XU444 n26 n1622 NETTRAN_DUMMY_3023 NETTRAN_DUMMY_3024 INV_X1 
XU443 n596 n1824 NETTRAN_DUMMY_3025 NETTRAN_DUMMY_3026 INV_X1 
XU442 n575 n1763 NETTRAN_DUMMY_3027 NETTRAN_DUMMY_3028 INV_X1 
XU441 n19 n1614 NETTRAN_DUMMY_3029 NETTRAN_DUMMY_3030 INV_X1 
XU440 n566 n1795 NETTRAN_DUMMY_3031 NETTRAN_DUMMY_3032 INV_X1 
XU437 n572 n1796 NETTRAN_DUMMY_3033 NETTRAN_DUMMY_3034 INV_X1 
XU419 n598 n1850 NETTRAN_DUMMY_3035 NETTRAN_DUMMY_3036 INV_X1 
XU418 n584 n1741 NETTRAN_DUMMY_3037 NETTRAN_DUMMY_3038 INV_X1 
XU417 n522 n1770 NETTRAN_DUMMY_3039 NETTRAN_DUMMY_3040 INV_X1 
XU416 n1531 n4 n248 n247 NETTRAN_DUMMY_3041 NETTRAN_DUMMY_3042 AND3_X1 
XU415 n625 n1758 NETTRAN_DUMMY_3043 NETTRAN_DUMMY_3044 INV_X1 
XU414 n1522 n1528 n410 NETTRAN_DUMMY_3045 NETTRAN_DUMMY_3046 NOR2_X1 
XU413 n606 n1779 NETTRAN_DUMMY_3047 NETTRAN_DUMMY_3048 INV_X1 
XU412 n204 n1650 NETTRAN_DUMMY_3049 NETTRAN_DUMMY_3050 INV_X1 
XU411 n541 n1767 NETTRAN_DUMMY_3051 NETTRAN_DUMMY_3052 INV_X1 
XU410 n553 n1674 NETTRAN_DUMMY_3053 NETTRAN_DUMMY_3054 INV_X1 
XU409 n31 n1625 NETTRAN_DUMMY_3055 NETTRAN_DUMMY_3056 INV_X1 
XU408 n603 n1759 NETTRAN_DUMMY_3057 NETTRAN_DUMMY_3058 INV_X1 
XU403 n605 n1778 NETTRAN_DUMMY_3059 NETTRAN_DUMMY_3060 INV_X1 
XU381 n4 n1610 NETTRAN_DUMMY_3061 NETTRAN_DUMMY_3062 INV_X1 
XU359 n626 n1844 NETTRAN_DUMMY_3063 NETTRAN_DUMMY_3064 INV_X1 
XU355 n547 n1833 NETTRAN_DUMMY_3065 NETTRAN_DUMMY_3066 INV_X1 
XU352 n564 n1775 NETTRAN_DUMMY_3067 NETTRAN_DUMMY_3068 INV_X1 
XU348 n620 n1841 NETTRAN_DUMMY_3069 NETTRAN_DUMMY_3070 INV_X1 
XU344 n530 n1771 NETTRAN_DUMMY_3071 NETTRAN_DUMMY_3072 INV_X1 
XU329 n550 n1790 NETTRAN_DUMMY_3073 NETTRAN_DUMMY_3074 INV_X1 
XU318 n10 n1646 NETTRAN_DUMMY_3075 NETTRAN_DUMMY_3076 INV_X1 
XU313 n585 n1742 NETTRAN_DUMMY_3077 NETTRAN_DUMMY_3078 INV_X1 
XU309 n560 n1808 NETTRAN_DUMMY_3079 NETTRAN_DUMMY_3080 INV_X1 
XU300 n557 n1789 NETTRAN_DUMMY_3081 NETTRAN_DUMMY_3082 INV_X1 
XU268 n527 n1811 NETTRAN_DUMMY_3083 NETTRAN_DUMMY_3084 INV_X1 
XU262 n578 n1832 NETTRAN_DUMMY_3085 NETTRAN_DUMMY_3086 INV_X1 
XU261 n559 n1765 NETTRAN_DUMMY_3087 NETTRAN_DUMMY_3088 INV_X1 
XU252 n587 n1743 NETTRAN_DUMMY_3089 NETTRAN_DUMMY_3090 INV_X1 
XU248 n619 n1826 NETTRAN_DUMMY_3091 NETTRAN_DUMMY_3092 INV_X1 
XU223 n588 n1805 NETTRAN_DUMMY_3093 NETTRAN_DUMMY_3094 INV_X1 
XU213 n571 n1776 NETTRAN_DUMMY_3095 NETTRAN_DUMMY_3096 INV_X1 
XU208 n552 n1754 NETTRAN_DUMMY_3097 NETTRAN_DUMMY_3098 INV_X1 
XU206 n589 n1797 NETTRAN_DUMMY_3099 NETTRAN_DUMMY_3100 INV_X1 
XU205 n532 n1791 NETTRAN_DUMMY_3101 NETTRAN_DUMMY_3102 INV_X1 
XU203 n590 n1761 NETTRAN_DUMMY_3103 NETTRAN_DUMMY_3104 INV_X1 
XU196 n609 n1745 NETTRAN_DUMMY_3105 NETTRAN_DUMMY_3106 INV_X1 
XU192 n497 n529 n742 NETTRAN_DUMMY_3107 NETTRAN_DUMMY_3108 NAND2_X1 
XU191 n502 n1745 n1230 NETTRAN_DUMMY_3109 NETTRAN_DUMMY_3110 NAND2_X1 
XU170 n1708 n1856 NETTRAN_DUMMY_3111 NETTRAN_DUMMY_3112 INV_X1 
XU168 n58 n1643 NETTRAN_DUMMY_3113 NETTRAN_DUMMY_3114 INV_X1 
XU130 n2 n4 n261 NETTRAN_DUMMY_3115 NETTRAN_DUMMY_3116 NAND2_X1 
XU106 n6 n10 n15 NETTRAN_DUMMY_3117 NETTRAN_DUMMY_3118 NAND2_X1 
XU58 addr[5] n451 NETTRAN_DUMMY_3119 NETTRAN_DUMMY_3120 INV_X1 
XU56 n448 n449 NETTRAN_DUMMY_3121 NETTRAN_DUMMY_3122 INV_X1 
XU55 n6 n4 n48 NETTRAN_DUMMY_3123 NETTRAN_DUMMY_3124 NAND2_X1 
XU53 n609 n502 n587 n1337 NETTRAN_DUMMY_3125 NETTRAN_DUMMY_3126 AOI21_X1 
XU44 n443 n444 NETTRAN_DUMMY_3127 NETTRAN_DUMMY_3128 INV_X1 
XU39 n7 n2 n27 NETTRAN_DUMMY_3129 NETTRAN_DUMMY_3130 NAND2_X1 
XU37 n519 n1522 n538 NETTRAN_DUMMY_3131 NETTRAN_DUMMY_3132 NAND2_X1 
XU30 n519 n520 n518 NETTRAN_DUMMY_3133 NETTRAN_DUMMY_3134 NAND2_X1 
XU22 n543 n1522 n558 NETTRAN_DUMMY_3135 NETTRAN_DUMMY_3136 NAND2_X1 
XU20 n497 n1701 n1694 NETTRAN_DUMMY_3137 NETTRAN_DUMMY_3138 NAND2_X1 
XU18 n520 n543 n542 NETTRAN_DUMMY_3139 NETTRAN_DUMMY_3140 NAND2_X1 
XU13 n9 n10 n8 NETTRAN_DUMMY_3141 NETTRAN_DUMMY_3142 NAND2_X1 
XU11 addr[7] n437 NETTRAN_DUMMY_3143 NETTRAN_DUMMY_3144 INV_X1 
XU9 n27 n1607 NETTRAN_DUMMY_3145 NETTRAN_DUMMY_3146 INV_X1 
XU8 n538 n1755 NETTRAN_DUMMY_3147 NETTRAN_DUMMY_3148 INV_X1 
XU7 n48 n1611 NETTRAN_DUMMY_3149 NETTRAN_DUMMY_3150 INV_X1 
XU6 n558 n1773 NETTRAN_DUMMY_3151 NETTRAN_DUMMY_3152 INV_X1 
XU5 n518 n1756 NETTRAN_DUMMY_3153 NETTRAN_DUMMY_3154 INV_X1 
XU4 n1688 n408 NETTRAN_DUMMY_3155 NETTRAN_DUMMY_3156 INV_X1 
XU3 n1664 n408 n409 NETTRAN_DUMMY_3157 NETTRAN_DUMMY_3158 NAND2_X1 
Xc1_reg_17_ n2059 clk_cts_0 n2022 NETTRAN_DUMMY_3159 NETTRAN_DUMMY_3160 NETTRAN_DUMMY_3161 DFF_X1 
XU1564 n629 n593 n462 n1519 NETTRAN_DUMMY_3162 NETTRAN_DUMMY_3163 MUX2_X1 
XU1563 n520 n528 n502 n1366 NETTRAN_DUMMY_3164 NETTRAN_DUMMY_3165 MUX2_X1 
XU1562 n1763 n1804 n502 n1354 NETTRAN_DUMMY_3166 NETTRAN_DUMMY_3167 MUX2_X1 
XU1561 n488 n517 n509 n1518 NETTRAN_DUMMY_3168 NETTRAN_DUMMY_3169 MUX2_X1 
XU1560 n1538 n1758 n502 n1517 NETTRAN_DUMMY_3170 NETTRAN_DUMMY_3171 MUX2_X1 
XU1559 n492 n1318 n509 n1516 NETTRAN_DUMMY_3172 NETTRAN_DUMMY_3173 MUX2_X1 
XU1558 n1505 n1765 n495 n1160 NETTRAN_DUMMY_3174 NETTRAN_DUMMY_3175 MUX2_X1 
XU543 addr[5] n1540 n46 NETTRAN_DUMMY_3176 NETTRAN_DUMMY_3177 NAND2_X1 
XU542 n1684 n1589 NETTRAN_DUMMY_3178 NETTRAN_DUMMY_3179 INV_X1 
XU541 n473 n1521 n750 NETTRAN_DUMMY_3180 NETTRAN_DUMMY_3181 NAND2_X1 
XU540 n1531 n448 n13 NETTRAN_DUMMY_3182 NETTRAN_DUMMY_3183 OR2_X1 
XU539 n4 n5 n3 NETTRAN_DUMMY_3184 NETTRAN_DUMMY_3185 NAND2_X1 
XU538 n531 n528 n582 NETTRAN_DUMMY_3186 NETTRAN_DUMMY_3187 NAND2_X1 
XU537 addr[7] n55 n248 NETTRAN_DUMMY_3188 NETTRAN_DUMMY_3189 NAND2_X1 
XU536 n464 n558 n1295 NETTRAN_DUMMY_3190 NETTRAN_DUMMY_3191 NAND2_X1 
XU535 n526 n543 n776 NETTRAN_DUMMY_3192 NETTRAN_DUMMY_3193 NAND2_X1 
XU533 addr[5] n2 n58 NETTRAN_DUMMY_3194 NETTRAN_DUMMY_3195 NAND2_X1 
XU531 n519 n526 n760 NETTRAN_DUMMY_3196 NETTRAN_DUMMY_3197 NAND2_X1 
XU530 n1701 n1702 n1690 NETTRAN_DUMMY_3198 NETTRAN_DUMMY_3199 NAND2_X1 
XU529 n448 n1537 n21 NETTRAN_DUMMY_3200 NETTRAN_DUMMY_3201 NAND2_X1 
XU528 n528 n519 n552 NETTRAN_DUMMY_3202 NETTRAN_DUMMY_3203 NAND2_X1 
XU527 n509 n1525 n587 NETTRAN_DUMMY_3204 NETTRAN_DUMMY_3205 NAND2_X1 
XU526 addr[5] n1531 n7 NETTRAN_DUMMY_3206 NETTRAN_DUMMY_3207 NAND2_X1 
XU525 n522 n528 n530 NETTRAN_DUMMY_3208 NETTRAN_DUMMY_3209 NAND2_X1 
XU524 addr[5] n1527 n130 NETTRAN_DUMMY_3210 NETTRAN_DUMMY_3211 NAND2_X1 
XU523 n513 n480 n524 NETTRAN_DUMMY_3212 NETTRAN_DUMMY_3213 NAND2_X1 
XU522 n6 n448 n19 NETTRAN_DUMMY_3214 NETTRAN_DUMMY_3215 NAND2_X1 
XU520 n501 IN0 n1685 NETTRAN_DUMMY_3216 NETTRAN_DUMMY_3217 NOR2_X1 
XU519 n531 n526 n560 NETTRAN_DUMMY_3218 NETTRAN_DUMMY_3219 NAND2_X1 
XU518 n517 n525 n545 NETTRAN_DUMMY_3220 NETTRAN_DUMMY_3221 NAND2_X1 
XU517 n517 n531 n541 NETTRAN_DUMMY_3222 NETTRAN_DUMMY_3223 NAND2_X1 
XU516 n515 n1526 n537 NETTRAN_DUMMY_3224 NETTRAN_DUMMY_3225 NAND2_X1 
XU515 n480 n513 n1726 NETTRAN_DUMMY_3226 NETTRAN_DUMMY_3227 NOR2_X1 
XU514 n480 n481 n1693 NETTRAN_DUMMY_3228 NETTRAN_DUMMY_3229 NOR2_X1 
XU512 n543 n517 n625 NETTRAN_DUMMY_3230 NETTRAN_DUMMY_3231 NAND2_X1 
XU511 n480 n1524 n1700 NETTRAN_DUMMY_3232 NETTRAN_DUMMY_3233 NOR2_X1 
XU510 n1589 n1700 n1701 n1676 NETTRAN_DUMMY_3234 NETTRAN_DUMMY_3235 OAI21_X1 
XU509 n528 n525 n527 NETTRAN_DUMMY_3236 NETTRAN_DUMMY_3237 NAND2_X1 
XU508 n448 n5 n10 NETTRAN_DUMMY_3238 NETTRAN_DUMMY_3239 NAND2_X1 
XU507 n521 n520 n548 NETTRAN_DUMMY_3240 NETTRAN_DUMMY_3241 NAND2_X1 
XU506 n5 n448 n411 NETTRAN_DUMMY_3242 NETTRAN_DUMMY_3243 XNOR2_X1 
XU505 n517 n522 n523 NETTRAN_DUMMY_3244 NETTRAN_DUMMY_3245 NAND2_X1 
XU503 n448 n486 n1680 NETTRAN_DUMMY_3246 NETTRAN_DUMMY_3247 NAND2_X1 
XU502 n513 n1318 n529 NETTRAN_DUMMY_3248 NETTRAN_DUMMY_3249 NAND2_X1 
XU501 n509 n1522 n522 NETTRAN_DUMMY_3250 NETTRAN_DUMMY_3251 NAND2_X1 
XU500 n448 n1 n4 NETTRAN_DUMMY_3252 NETTRAN_DUMMY_3253 NAND2_X1 
XU499 n509 n528 n543 NETTRAN_DUMMY_3254 NETTRAN_DUMMY_3255 NAND2_X1 
XU496 IN0 n501 n1708 NETTRAN_DUMMY_3256 NETTRAN_DUMMY_3257 NAND2_X1 
XU495 n509 n517 n519 NETTRAN_DUMMY_3258 NETTRAN_DUMMY_3259 NAND2_X1 
XU493 n509 n520 n531 NETTRAN_DUMMY_3260 NETTRAN_DUMMY_3261 NAND2_X1 
XU492 n513 n497 n6 NETTRAN_DUMMY_3262 NETTRAN_DUMMY_3263 NAND2_X1 
XU490 n533 n525 n532 NETTRAN_DUMMY_3264 NETTRAN_DUMMY_3265 NAND2_X1 
XU489 n509 n526 n525 NETTRAN_DUMMY_3266 NETTRAN_DUMMY_3267 NAND2_X1 
XU488 n480 IN0 n1701 NETTRAN_DUMMY_3268 NETTRAN_DUMMY_3269 NOR2_X1 
XU487 n460 n461 NETTRAN_DUMMY_3270 NETTRAN_DUMMY_3271 INV_X1 
XU482 addr[0] n501 n2 NETTRAN_DUMMY_3272 NETTRAN_DUMMY_3273 NAND2_X1 
XU480 n492 n480 n520 NETTRAN_DUMMY_3274 NETTRAN_DUMMY_3275 NAND2_X1 
XU479 n1680 n1664 NETTRAN_DUMMY_3276 NETTRAN_DUMMY_3277 INV_X1 
XU478 n39 n1630 NETTRAN_DUMMY_3278 NETTRAN_DUMMY_3279 INV_X1 
XU477 n18 n1613 NETTRAN_DUMMY_3280 NETTRAN_DUMMY_3281 INV_X1 
XU476 n1517 n1757 NETTRAN_DUMMY_3282 NETTRAN_DUMMY_3283 INV_X1 
XU475 n1300 n519 n1307 NETTRAN_DUMMY_3284 NETTRAN_DUMMY_3285 AND2_X1 
XU474 n607 n1840 NETTRAN_DUMMY_3286 NETTRAN_DUMMY_3287 INV_X1 
XU473 n34 n1628 NETTRAN_DUMMY_3288 NETTRAN_DUMMY_3289 INV_X1 
XU472 n24 n1620 NETTRAN_DUMMY_3290 NETTRAN_DUMMY_3291 INV_X1 
XU471 n50 n1639 NETTRAN_DUMMY_3292 NETTRAN_DUMMY_3293 INV_X1 
XU470 n47 n1637 NETTRAN_DUMMY_3294 NETTRAN_DUMMY_3295 INV_X1 
XU469 n20 n1616 NETTRAN_DUMMY_3296 NETTRAN_DUMMY_3297 INV_X1 
XU468 n221 n1645 NETTRAN_DUMMY_3298 NETTRAN_DUMMY_3299 INV_X1 
XU467 n613 n1845 NETTRAN_DUMMY_3300 NETTRAN_DUMMY_3301 INV_X1 
XU466 n3 n1612 NETTRAN_DUMMY_3302 NETTRAN_DUMMY_3303 INV_X1 
XU465 n611 n1831 NETTRAN_DUMMY_3304 NETTRAN_DUMMY_3305 INV_X1 
XU464 n610 n1784 NETTRAN_DUMMY_3306 NETTRAN_DUMMY_3307 INV_X1 
XU463 n56 n1641 NETTRAN_DUMMY_3308 NETTRAN_DUMMY_3309 INV_X1 
XU462 n32 n1626 NETTRAN_DUMMY_3310 NETTRAN_DUMMY_3311 INV_X1 
XU461 n22 n1618 NETTRAN_DUMMY_3312 NETTRAN_DUMMY_3313 INV_X1 
XU460 n591 n1777 NETTRAN_DUMMY_3314 NETTRAN_DUMMY_3315 INV_X1 
XU459 n595 n1804 NETTRAN_DUMMY_3316 NETTRAN_DUMMY_3317 INV_X1 
XU458 n570 n1846 NETTRAN_DUMMY_3318 NETTRAN_DUMMY_3319 INV_X1 
XU457 n1633 n248 n354 NETTRAN_DUMMY_3320 NETTRAN_DUMMY_3321 NAND2_X1 
XU456 n542 n1836 NETTRAN_DUMMY_3322 NETTRAN_DUMMY_3323 INV_X1 
XU455 n1836 n1295 n1294 NETTRAN_DUMMY_3324 NETTRAN_DUMMY_3325 NAND2_X1 
XU454 n51 n1640 NETTRAN_DUMMY_3326 NETTRAN_DUMMY_3327 INV_X1 
XU453 n582 n1838 NETTRAN_DUMMY_3328 NETTRAN_DUMMY_3329 INV_X1 
XU452 n49 n1638 NETTRAN_DUMMY_3330 NETTRAN_DUMMY_3331 INV_X1 
XU451 n576 n1839 NETTRAN_DUMMY_3332 NETTRAN_DUMMY_3333 INV_X1 
XU1162 n519 n1753 NETTRAN_DUMMY_3334 NETTRAN_DUMMY_3335 INV_X1 
XU1158 n513 n501 n736 NETTRAN_DUMMY_3336 NETTRAN_DUMMY_3337 NAND2_X1 
XU1156 n1188 n1186 n1200 NETTRAN_DUMMY_3338 NETTRAN_DUMMY_3339 NOR2_X1 
XU1152 n220 n223 addr[3] n222 NETTRAN_DUMMY_3340 NETTRAN_DUMMY_3341 AOI21_X1 
XU1134 n578 n501 n1086 NETTRAN_DUMMY_3342 NETTRAN_DUMMY_3343 AND2_X1 
XU1131 n443 n517 n844 NETTRAN_DUMMY_3344 NETTRAN_DUMMY_3345 NOR2_X1 
XU1129 n442 n1547 n638 NETTRAN_DUMMY_3346 NETTRAN_DUMMY_3347 NOR2_X1 
XU1112 IN0 n1650 n168 NETTRAN_DUMMY_3348 NETTRAN_DUMMY_3349 NOR2_X1 
XU1104 n585 n507 n627 n1406 NETTRAN_DUMMY_3350 NETTRAN_DUMMY_3351 AOI21_X1 
XU1102 n1752 n453 n536 n1286 NETTRAN_DUMMY_3352 NETTRAN_DUMMY_3353 AOI21_X1 
XU1080 n593 n501 n579 n932 NETTRAN_DUMMY_3354 NETTRAN_DUMMY_3355 OAI21_X1 
XU1074 n608 n1785 NETTRAN_DUMMY_3356 NETTRAN_DUMMY_3357 INV_X1 
XU1045 n443 n1790 n794 NETTRAN_DUMMY_3358 NETTRAN_DUMMY_3359 NOR2_X1 
XU1043 n59 n1642 NETTRAN_DUMMY_3360 NETTRAN_DUMMY_3361 INV_X1 
XU1015 n57 n1644 NETTRAN_DUMMY_3362 NETTRAN_DUMMY_3363 INV_X1 
XU1012 n13 n1608 NETTRAN_DUMMY_3364 NETTRAN_DUMMY_3365 INV_X1 
XU1011 n407 n1603 NETTRAN_DUMMY_3366 NETTRAN_DUMMY_3367 INV_X1 
XU986 n17 n1609 NETTRAN_DUMMY_3368 NETTRAN_DUMMY_3369 INV_X1 
XU984 n25 n1621 NETTRAN_DUMMY_3370 NETTRAN_DUMMY_3371 INV_X1 
XU956 n540 n1847 NETTRAN_DUMMY_3372 NETTRAN_DUMMY_3373 INV_X1 
XU947 n817 n1781 NETTRAN_DUMMY_3374 NETTRAN_DUMMY_3375 INV_X1 
XU927 n468 n1539 n692 NETTRAN_DUMMY_3376 NETTRAN_DUMMY_3377 NOR2_X1 
XU925 n452 n534 n694 NETTRAN_DUMMY_3378 NETTRAN_DUMMY_3379 NOR2_X1 
XU911 n473 n965 n969 NETTRAN_DUMMY_3380 NETTRAN_DUMMY_3381 NOR2_X1 
XU898 n462 n936 n940 NETTRAN_DUMMY_3382 NETTRAN_DUMMY_3383 NOR2_X1 
XU887 n521 n526 n1369 NETTRAN_DUMMY_3384 NETTRAN_DUMMY_3385 NAND2_X1 
XU883 n341 n347 n433 n346 NETTRAN_DUMMY_3386 NETTRAN_DUMMY_3387 AOI21_X1 
XU869 n1643 n460 n13 n379 NETTRAN_DUMMY_3388 NETTRAN_DUMMY_3389 AOI21_X1 
XU858 n11 n1591 NETTRAN_DUMMY_3390 NETTRAN_DUMMY_3391 INV_X1 
XU851 n535 n1295 n1448 NETTRAN_DUMMY_3392 NETTRAN_DUMMY_3393 NAND2_X1 
XU840 n1116 n1108 n1109 n1115 NETTRAN_DUMMY_3394 NETTRAN_DUMMY_3395 OAI21_X1 
XU838 n42 n1633 NETTRAN_DUMMY_3396 NETTRAN_DUMMY_3397 INV_X1 
XU831 n604 n1853 NETTRAN_DUMMY_3398 NETTRAN_DUMMY_3399 INV_X1 
XU811 n29 n1594 NETTRAN_DUMMY_3400 NETTRAN_DUMMY_3401 INV_X1 
XU809 n554 n1772 NETTRAN_DUMMY_3402 NETTRAN_DUMMY_3403 INV_X1 
XU790 n501 n569 n743 NETTRAN_DUMMY_3404 NETTRAN_DUMMY_3405 NOR2_X1 
XU779 n555 n1855 NETTRAN_DUMMY_3406 NETTRAN_DUMMY_3407 INV_X1 
XU775 n586 n1762 NETTRAN_DUMMY_3408 NETTRAN_DUMMY_3409 INV_X1 
XU765 n445 n448 n1687 n1706 NETTRAN_DUMMY_3410 NETTRAN_DUMMY_3411 OAI21_X1 
XU757 n1706 n1590 NETTRAN_DUMMY_3412 NETTRAN_DUMMY_3413 INV_X1 
XU756 n38 n1597 NETTRAN_DUMMY_3414 NETTRAN_DUMMY_3415 INV_X1 
XU754 n35 n1595 NETTRAN_DUMMY_3416 NETTRAN_DUMMY_3417 INV_X1 
XU750 n41 n1632 NETTRAN_DUMMY_3418 NETTRAN_DUMMY_3419 INV_X1 
XU748 n8 n1648 NETTRAN_DUMMY_3420 NETTRAN_DUMMY_3421 INV_X1 
XU747 n402 n403 n401 NETTRAN_DUMMY_3422 NETTRAN_DUMMY_3423 NAND2_X1 
XU731 n1661 n487 n23 n298 NETTRAN_DUMMY_3424 NETTRAN_DUMMY_3425 AOI21_X1 
XU728 n55 n1600 NETTRAN_DUMMY_3426 NETTRAN_DUMMY_3427 INV_X1 
XU726 n1599 n484 n311 n310 NETTRAN_DUMMY_3428 NETTRAN_DUMMY_3429 AOI21_X1 
XU724 n581 n1849 NETTRAN_DUMMY_3430 NETTRAN_DUMMY_3431 INV_X1 
XU705 n524 n1849 n501 n1325 NETTRAN_DUMMY_3432 NETTRAN_DUMMY_3433 OAI21_X1 
XU702 n1510 n1752 NETTRAN_DUMMY_3434 NETTRAN_DUMMY_3435 INV_X1 
XU687 n416 n1654 NETTRAN_DUMMY_3436 NETTRAN_DUMMY_3437 INV_X1 
XU677 n44 n1635 NETTRAN_DUMMY_3438 NETTRAN_DUMMY_3439 INV_X1 
XU671 n415 n1653 NETTRAN_DUMMY_3440 NETTRAN_DUMMY_3441 INV_X1 
XU649 n419 n1656 NETTRAN_DUMMY_3442 NETTRAN_DUMMY_3443 INV_X1 
XU646 n418 n1655 NETTRAN_DUMMY_3444 NETTRAN_DUMMY_3445 INV_X1 
XU636 n414 n1652 NETTRAN_DUMMY_3446 NETTRAN_DUMMY_3447 INV_X1 
XU635 n1502 n1663 NETTRAN_DUMMY_3448 NETTRAN_DUMMY_3449 INV_X1 
XU627 n1519 n1673 NETTRAN_DUMMY_3450 NETTRAN_DUMMY_3451 INV_X1 
XU618 n422 n1659 NETTRAN_DUMMY_3452 NETTRAN_DUMMY_3453 INV_X1 
XU615 n1511 n1672 NETTRAN_DUMMY_3454 NETTRAN_DUMMY_3455 INV_X1 
XU611 n1520 n509 n607 NETTRAN_DUMMY_3456 NETTRAN_DUMMY_3457 NAND2_X1 
XU608 n473 n1499 n1110 NETTRAN_DUMMY_3458 NETTRAN_DUMMY_3459 NAND2_X1 
XU604 addr[7] n28 n351 NETTRAN_DUMMY_3460 NETTRAN_DUMMY_3461 NOR2_X1 
XU603 n433 n522 n993 NETTRAN_DUMMY_3462 NETTRAN_DUMMY_3463 NOR2_X1 
XU598 n442 n1539 n710 NETTRAN_DUMMY_3464 NETTRAN_DUMMY_3465 NOR2_X1 
XU593 n480 n1524 n198 NETTRAN_DUMMY_3466 NETTRAN_DUMMY_3467 NOR2_X1 
XU592 n462 n1051 n1055 NETTRAN_DUMMY_3468 NETTRAN_DUMMY_3469 NOR2_X1 
XU591 n417 n1598 NETTRAN_DUMMY_3470 NETTRAN_DUMMY_3471 INV_X1 
XU579 n1 n19 n54 NETTRAN_DUMMY_3472 NETTRAN_DUMMY_3473 NAND2_X1 
XU570 n616 n1783 NETTRAN_DUMMY_3474 NETTRAN_DUMMY_3475 INV_X1 
XU565 n579 n1812 NETTRAN_DUMMY_3476 NETTRAN_DUMMY_3477 INV_X1 
XU562 n1524 addr[5] n43 NETTRAN_DUMMY_3478 NETTRAN_DUMMY_3479 NAND2_X1 
XU561 n1743 n502 n561 n1166 NETTRAN_DUMMY_3480 NETTRAN_DUMMY_3481 AOI21_X1 
XU560 n1765 n473 n527 n869 NETTRAN_DUMMY_3482 NETTRAN_DUMMY_3483 AOI21_X1 
XU559 n1816 n477 n571 n1024 NETTRAN_DUMMY_3484 NETTRAN_DUMMY_3485 AOI21_X1 
XU558 n5 n19 n105 NETTRAN_DUMMY_3486 NETTRAN_DUMMY_3487 NAND2_X1 
XU555 n471 n472 NETTRAN_DUMMY_3488 NETTRAN_DUMMY_3489 INV_X1 
XU553 n54 n1615 NETTRAN_DUMMY_3490 NETTRAN_DUMMY_3491 INV_X1 
XU552 n17 addr[7] n53 n252 NETTRAN_DUMMY_3492 NETTRAN_DUMMY_3493 AOI21_X1 
XU551 n501 n448 n204 NETTRAN_DUMMY_3494 NETTRAN_DUMMY_3495 NAND2_X1 
XU550 n1543 n453 n565 n1276 NETTRAN_DUMMY_3496 NETTRAN_DUMMY_3497 AOI21_X1 
XU549 n1586 n1690 n468 n1689 NETTRAN_DUMMY_3498 NETTRAN_DUMMY_3499 NAND3_X1 
XU548 n1689 n1687 n1688 n1678 NETTRAN_DUMMY_3500 NETTRAN_DUMMY_3501 OAI21_X1 
XU547 n464 n563 n1300 NETTRAN_DUMMY_3502 NETTRAN_DUMMY_3503 NAND2_X1 
XU546 n561 n1774 NETTRAN_DUMMY_3504 NETTRAN_DUMMY_3505 INV_X1 
XU545 n58 n5 n57 NETTRAN_DUMMY_3506 NETTRAN_DUMMY_3507 NAND2_X1 
XU544 n1523 n502 n616 n1204 NETTRAN_DUMMY_3508 NETTRAN_DUMMY_3509 AOI21_X1 
XU1616 n492 n493 NETTRAN_DUMMY_3510 NETTRAN_DUMMY_3511 INV_X1 
XU1614 n480 n493 n528 NETTRAN_DUMMY_3512 NETTRAN_DUMMY_3513 NAND2_X1 
XU1613 n488 n493 n526 NETTRAN_DUMMY_3514 NETTRAN_DUMMY_3515 NAND2_X1 
XU1612 n492 n488 n517 NETTRAN_DUMMY_3516 NETTRAN_DUMMY_3517 NAND2_X1 
XU1611 n624 n1666 NETTRAN_DUMMY_3518 NETTRAN_DUMMY_3519 INV_X1 
XU1610 n452 n1666 n1187 NETTRAN_DUMMY_3520 NETTRAN_DUMMY_3521 NAND2_X1 
XU1609 n1697 addr[0] n1728 NETTRAN_DUMMY_3522 NETTRAN_DUMMY_3523 AND2_X1 
XU1608 n52 n1599 NETTRAN_DUMMY_3524 NETTRAN_DUMMY_3525 INV_X1 
XU1607 n484 n1536 n189 NETTRAN_DUMMY_3526 NETTRAN_DUMMY_3527 NAND2_X1 
XU1606 n1704 n1586 NETTRAN_DUMMY_3528 NETTRAN_DUMMY_3529 INV_X1 
XU1605 n1680 n1704 n1697 NETTRAN_DUMMY_3530 NETTRAN_DUMMY_3531 NOR2_X1 
XU1603 n433 n442 n1688 NETTRAN_DUMMY_3532 NETTRAN_DUMMY_3533 NAND2_X1 
XU1602 n487 n486 n1682 NETTRAN_DUMMY_3534 NETTRAN_DUMMY_3535 NAND2_X1 
XU1601 n1684 n442 IN0 n1729 NETTRAN_DUMMY_3536 NETTRAN_DUMMY_3537 OAI21_X1 
XU1600 n448 n442 n1699 NETTRAN_DUMMY_3538 NETTRAN_DUMMY_3539 NOR2_X1 
XU1598 n487 n488 NETTRAN_DUMMY_3540 NETTRAN_DUMMY_3541 INV_X2 
XU1589 n30 n1624 NETTRAN_DUMMY_3542 NETTRAN_DUMMY_3543 INV_X1 
XU1588 n46 n1636 NETTRAN_DUMMY_3544 NETTRAN_DUMMY_3545 INV_X1 
XU1587 n1508 n1806 NETTRAN_DUMMY_3546 NETTRAN_DUMMY_3547 INV_X1 
XU1586 n1512 n1749 NETTRAN_DUMMY_3548 NETTRAN_DUMMY_3549 INV_X1 
XU1585 n420 n1657 NETTRAN_DUMMY_3550 NETTRAN_DUMMY_3551 INV_X1 
XU1584 n1516 n1828 NETTRAN_DUMMY_3552 NETTRAN_DUMMY_3553 INV_X1 
XU1583 n1503 n1670 NETTRAN_DUMMY_3554 NETTRAN_DUMMY_3555 INV_X1 
XU1582 n28 n1623 NETTRAN_DUMMY_3556 NETTRAN_DUMMY_3557 INV_X1 
XU1581 n412 n1604 NETTRAN_DUMMY_3558 NETTRAN_DUMMY_3559 INV_X1 
XU1580 n423 n1660 NETTRAN_DUMMY_3560 NETTRAN_DUMMY_3561 INV_X1 
XU1579 n421 n1658 NETTRAN_DUMMY_3562 NETTRAN_DUMMY_3563 INV_X1 
XU1578 n425 n1662 NETTRAN_DUMMY_3564 NETTRAN_DUMMY_3565 INV_X1 
XU1577 n1300 n837 n1299 NETTRAN_DUMMY_3566 NETTRAN_DUMMY_3567 AND2_X1 
XU1576 n37 n1629 NETTRAN_DUMMY_3568 NETTRAN_DUMMY_3569 INV_X1 
XU1575 n1505 n1817 NETTRAN_DUMMY_3570 NETTRAN_DUMMY_3571 INV_X1 
XU1574 n549 n1822 NETTRAN_DUMMY_3572 NETTRAN_DUMMY_3573 INV_X1 
XU1573 n521 n1768 NETTRAN_DUMMY_3574 NETTRAN_DUMMY_3575 INV_X1 
XU1572 n1498 n1668 NETTRAN_DUMMY_3576 NETTRAN_DUMMY_3577 INV_X1 
XU1571 n484 n430 n1540 n317 NETTRAN_DUMMY_3578 NETTRAN_DUMMY_3579 OAI21_X1 
XU1570 n1635 n317 n316 NETTRAN_DUMMY_3580 NETTRAN_DUMMY_3581 NAND2_X1 
XU1569 n130 n1649 NETTRAN_DUMMY_3582 NETTRAN_DUMMY_3583 INV_X1 
XU1568 n621 n1748 NETTRAN_DUMMY_3584 NETTRAN_DUMMY_3585 INV_X1 
XU1567 n618 n1747 NETTRAN_DUMMY_3586 NETTRAN_DUMMY_3587 INV_X1 
XU1566 n632 n1667 NETTRAN_DUMMY_3588 NETTRAN_DUMMY_3589 INV_X1 
XU1565 n615 n1780 NETTRAN_DUMMY_3590 NETTRAN_DUMMY_3591 INV_X1 
XU1555 n617 n1746 NETTRAN_DUMMY_3592 NETTRAN_DUMMY_3593 INV_X1 
XU1536 n40 n1631 NETTRAN_DUMMY_3594 NETTRAN_DUMMY_3595 INV_X1 
XU1535 n599 n1814 NETTRAN_DUMMY_3596 NETTRAN_DUMMY_3597 INV_X1 
XU1534 n424 n1661 NETTRAN_DUMMY_3598 NETTRAN_DUMMY_3599 INV_X1 
XU1533 n837 n1842 NETTRAN_DUMMY_3600 NETTRAN_DUMMY_3601 INV_X1 
XU1532 n602 n1815 NETTRAN_DUMMY_3602 NETTRAN_DUMMY_3603 INV_X1 
XU1531 n544 n1852 NETTRAN_DUMMY_3604 NETTRAN_DUMMY_3605 INV_X1 
XU1530 n614 n1825 NETTRAN_DUMMY_3606 NETTRAN_DUMMY_3607 INV_X1 
XU1529 n592 n1744 NETTRAN_DUMMY_3608 NETTRAN_DUMMY_3609 INV_X1 
XU1528 n573 n1787 NETTRAN_DUMMY_3610 NETTRAN_DUMMY_3611 INV_X1 
XU1527 n311 n1605 NETTRAN_DUMMY_3612 NETTRAN_DUMMY_3613 INV_X1 
XU1474 n36 n1596 NETTRAN_DUMMY_3614 NETTRAN_DUMMY_3615 INV_X1 
XU1454 n1685 n445 n1683 NETTRAN_DUMMY_3616 NETTRAN_DUMMY_3617 OR2_X1 
XU1436 n594 n1760 NETTRAN_DUMMY_3618 NETTRAN_DUMMY_3619 INV_X1 
XU1430 n33 n1627 NETTRAN_DUMMY_3620 NETTRAN_DUMMY_3621 INV_X1 
XU1392 n463 n731 n732 NETTRAN_DUMMY_3622 NETTRAN_DUMMY_3623 NOR2_X1 
XU1389 n734 n501 n733 NETTRAN_DUMMY_3624 NETTRAN_DUMMY_3625 NAND2_X1 
XU1378 n1366 n525 n1365 NETTRAN_DUMMY_3626 NETTRAN_DUMMY_3627 NAND2_X1 
XU1361 n525 n501 n589 n1171 NETTRAN_DUMMY_3628 NETTRAN_DUMMY_3629 OAI21_X1 
XU1349 n477 n588 n1411 NETTRAN_DUMMY_3630 NETTRAN_DUMMY_3631 NAND2_X1 
XU1346 n585 n501 n1322 NETTRAN_DUMMY_3632 NETTRAN_DUMMY_3633 AND2_X1 
XU1333 n626 n464 n529 n1310 NETTRAN_DUMMY_3634 NETTRAN_DUMMY_3635 AOI21_X1 
XU1330 n537 n501 n1229 NETTRAN_DUMMY_3636 NETTRAN_DUMMY_3637 NOR2_X1 
XU1323 n546 n1585 NETTRAN_DUMMY_3638 NETTRAN_DUMMY_3639 INV_X1 
XU1319 n462 n1543 n1094 NETTRAN_DUMMY_3640 NETTRAN_DUMMY_3641 NOR2_X1 
XU1316 n1853 n507 n910 NETTRAN_DUMMY_3642 NETTRAN_DUMMY_3643 NAND2_X1 
XU1310 n462 n908 n912 NETTRAN_DUMMY_3644 NETTRAN_DUMMY_3645 NOR2_X1 
XU1300 n445 n1541 n635 NETTRAN_DUMMY_3646 NETTRAN_DUMMY_3647 NOR2_X1 
XU1253 n562 n1848 NETTRAN_DUMMY_3648 NETTRAN_DUMMY_3649 INV_X1 
XU1252 n448 n1524 n342 NETTRAN_DUMMY_3650 NETTRAN_DUMMY_3651 NOR2_X1 
XU1228 n2 n10 n328 NETTRAN_DUMMY_3652 NETTRAN_DUMMY_3653 NAND2_X1 
XU1225 n15 n1647 NETTRAN_DUMMY_3654 NETTRAN_DUMMY_3655 INV_X1 
XU1220 n7 n1606 NETTRAN_DUMMY_3656 NETTRAN_DUMMY_3657 INV_X1 
XU1212 n23 n1619 NETTRAN_DUMMY_3658 NETTRAN_DUMMY_3659 INV_X1 
XU1210 n406 n1602 NETTRAN_DUMMY_3660 NETTRAN_DUMMY_3661 INV_X1 
XU1207 n435 n1744 n997 NETTRAN_DUMMY_3662 NETTRAN_DUMMY_3663 NOR2_X1 
XU1190 n600 n821 n825 NETTRAN_DUMMY_3664 NETTRAN_DUMMY_3665 NOR2_X1 
XU1185 n16 n1593 NETTRAN_DUMMY_3666 NETTRAN_DUMMY_3667 INV_X1 
XU1179 n1537 n1643 n358 NETTRAN_DUMMY_3668 NETTRAN_DUMMY_3669 NOR2_X1 
XU1711 n1524 n1729 n472 n434 n1717 NETTRAN_DUMMY_3670 NETTRAN_DUMMY_3671 NAND4_X1 
XU1710 n1586 n497 n448 n1713 n1716 NETTRAN_DUMMY_3672 NETTRAN_DUMMY_3673 OAI211_X1 
XU1709 n1716 n1717 n1718 n1719 N13521 NETTRAN_DUMMY_3674 NETTRAN_DUMMY_3675 NAND4_X1 
XU1708 n1522 n516 n521 NETTRAN_DUMMY_3676 NETTRAN_DUMMY_3677 OR2_X1 
XU1707 n513 n493 n1686 NETTRAN_DUMMY_3678 NETTRAN_DUMMY_3679 NOR2_X1 
XU1706 n488 n1686 n1856 n1681 NETTRAN_DUMMY_3680 NETTRAN_DUMMY_3681 OAI21_X1 
XU1705 n501 n516 n1702 NETTRAN_DUMMY_3682 NETTRAN_DUMMY_3683 NAND2_X1 
XU1704 n1520 n516 n837 NETTRAN_DUMMY_3684 NETTRAN_DUMMY_3685 NAND2_X1 
XU1703 n1693 n461 n1687 NETTRAN_DUMMY_3686 NETTRAN_DUMMY_3687 NAND2_X1 
XU1702 n5 n493 n45 NETTRAN_DUMMY_3688 NETTRAN_DUMMY_3689 NAND2_X1 
XU1701 n509 n493 n544 NETTRAN_DUMMY_3690 NETTRAN_DUMMY_3691 NAND2_X1 
XU1700 n577 n628 n444 n717 NETTRAN_DUMMY_3692 NETTRAN_DUMMY_3693 OAI21_X1 
XU1699 n461 n1762 n444 n600 NETTRAN_DUMMY_3694 NETTRAN_DUMMY_3695 AOI21_X1 
XU1698 n501 n488 addr[0] n1734 NETTRAN_DUMMY_3696 NETTRAN_DUMMY_3697 NAND3_X1 
XU1697 n468 n1694 n1734 n1732 NETTRAN_DUMMY_3698 NETTRAN_DUMMY_3699 AOI21_X1 
XU1696 n2 n451 n29 NETTRAN_DUMMY_3700 NETTRAN_DUMMY_3701 NAND2_X1 
XU1695 n1522 n516 n817 NETTRAN_DUMMY_3702 NETTRAN_DUMMY_3703 NAND2_X1 
XU1694 n444 n1690 n468 n1695 NETTRAN_DUMMY_3704 NETTRAN_DUMMY_3705 AOI21_X1 
XU1693 n1695 n1587 NETTRAN_DUMMY_3706 NETTRAN_DUMMY_3707 INV_X1 
XU1692 n1587 n468 n1685 n1691 NETTRAN_DUMMY_3708 NETTRAN_DUMMY_3709 OAI21_X1 
XU1691 n535 n472 n1528 n534 NETTRAN_DUMMY_3710 NETTRAN_DUMMY_3711 OAI21_X1 
XU1690 addr[0] n449 n311 NETTRAN_DUMMY_3712 NETTRAN_DUMMY_3713 NAND2_X1 
XU1689 n512 n517 n897 NETTRAN_DUMMY_3714 NETTRAN_DUMMY_3715 NAND2_X1 
XU1688 n520 n461 n574 NETTRAN_DUMMY_3716 NETTRAN_DUMMY_3717 NAND2_X1 
XU1687 n512 n433 n488 n1725 NETTRAN_DUMMY_3718 NETTRAN_DUMMY_3719 OAI21_X1 
XU1686 n1725 n501 n1726 n497 n1723 NETTRAN_DUMMY_3720 NETTRAN_DUMMY_3721 AOI22_X1 
XU1685 n1524 n451 n36 NETTRAN_DUMMY_3722 NETTRAN_DUMMY_3723 NAND2_X1 
XU1684 n488 n512 n551 NETTRAN_DUMMY_3724 NETTRAN_DUMMY_3725 NAND2_X1 
XU1683 n512 n528 n540 NETTRAN_DUMMY_3726 NETTRAN_DUMMY_3727 NAND2_X1 
XU1682 addr[1] n449 n38 NETTRAN_DUMMY_3728 NETTRAN_DUMMY_3729 NAND2_X1 
XU1681 n468 n1693 n472 n1694 n1692 NETTRAN_DUMMY_3730 NETTRAN_DUMMY_3731 OAI22_X1 
XU1680 n480 n512 n581 NETTRAN_DUMMY_3732 NETTRAN_DUMMY_3733 NAND2_X1 
XU1679 n512 n1526 n539 NETTRAN_DUMMY_3734 NETTRAN_DUMMY_3735 NAND2_X1 
XU1678 n1676 n1588 NETTRAN_DUMMY_3736 NETTRAN_DUMMY_3737 INV_X1 
XU1677 n1694 n486 n1698 NETTRAN_DUMMY_3738 NETTRAN_DUMMY_3739 AND2_X1 
XU1676 n1588 n1697 n1690 n1698 n1699 n1696 NETTRAN_DUMMY_3740 NETTRAN_DUMMY_3741 AOI221_X1 
XU1675 n1696 n1590 n434 n486 n1684 N4870 NETTRAN_DUMMY_3742 NETTRAN_DUMMY_3743 OAI221_X1 
XU1674 n1684 n1680 n1681 n1682 n1683 n1679 NETTRAN_DUMMY_3744 NETTRAN_DUMMY_3745 OAI221_X1 
XU1673 n448 n1691 n1692 n444 n1675 NETTRAN_DUMMY_3746 NETTRAN_DUMMY_3747 AOI22_X1 
XU1672 n1678 n449 n433 n1679 n1677 NETTRAN_DUMMY_3748 NETTRAN_DUMMY_3749 AOI22_X1 
XU1671 n1677 n433 n1675 n461 n1676 N5090 NETTRAN_DUMMY_3750 NETTRAN_DUMMY_3751 OAI221_X1 
XU1670 n501 n1726 n472 n1736 NETTRAN_DUMMY_3752 NETTRAN_DUMMY_3753 NOR3_X1 
XU1669 n1732 n1586 n1733 n1731 NETTRAN_DUMMY_3754 NETTRAN_DUMMY_3755 NOR3_X1 
XU1668 n1736 n1735 n461 n1730 NETTRAN_DUMMY_3756 NETTRAN_DUMMY_3757 AOI21_X1 
XU1667 n1731 n452 n1730 n1664 n434 N13331 NETTRAN_DUMMY_3758 NETTRAN_DUMMY_3759 OAI221_X1 
XU1666 n520 n512 n569 NETTRAN_DUMMY_3760 NETTRAN_DUMMY_3761 NAND2_X1 
XU1665 n1318 n512 n535 NETTRAN_DUMMY_3762 NETTRAN_DUMMY_3763 NAND2_X1 
XU1664 n445 n1680 n1701 n1715 NETTRAN_DUMMY_3764 NETTRAN_DUMMY_3765 OAI21_X1 
XU1663 addr[0] n1715 n1684 n1714 NETTRAN_DUMMY_3766 NETTRAN_DUMMY_3767 AOI21_X1 
XU1662 n1714 n1713 n1699 n472 n1589 n1712 NETTRAN_DUMMY_3768 NETTRAN_DUMMY_3769 AOI221_X1 
XU1661 n492 n512 n555 NETTRAN_DUMMY_3770 NETTRAN_DUMMY_3771 NAND2_X1 
XU1660 n513 n488 n593 NETTRAN_DUMMY_3772 NETTRAN_DUMMY_3773 NAND2_X1 
XU1659 n512 n526 n536 NETTRAN_DUMMY_3774 NETTRAN_DUMMY_3775 NAND2_X1 
XU1658 n526 n1526 NETTRAN_DUMMY_3776 NETTRAN_DUMMY_3777 INV_X1 
XU1657 n448 n444 n1684 NETTRAN_DUMMY_3778 NETTRAN_DUMMY_3779 NAND2_X1 
XU1656 n1724 n1722 n1708 n1723 n461 n1720 NETTRAN_DUMMY_3780 NETTRAN_DUMMY_3781 OAI221_X1 
XU1655 n434 n442 n1524 n1721 NETTRAN_DUMMY_3782 NETTRAN_DUMMY_3783 NOR3_X1 
XU1654 n1721 n408 n1680 n1699 n1720 n1719 NETTRAN_DUMMY_3784 NETTRAN_DUMMY_3785 AOI221_X1 
XU1653 n512 n497 n1 NETTRAN_DUMMY_3786 NETTRAN_DUMMY_3787 NAND2_X1 
XU1652 n533 n512 n616 NETTRAN_DUMMY_3788 NETTRAN_DUMMY_3789 NAND2_X1 
XU1651 n517 n1525 NETTRAN_DUMMY_3790 NETTRAN_DUMMY_3791 INV_X1 
XU1650 n501 n516 n5 NETTRAN_DUMMY_3792 NETTRAN_DUMMY_3793 NAND2_X1 
XU1649 n5 n1524 NETTRAN_DUMMY_3794 NETTRAN_DUMMY_3795 INV_X1 
XU1648 n583 n1523 NETTRAN_DUMMY_3796 NETTRAN_DUMMY_3797 INV_X1 
XU1647 n533 n1522 NETTRAN_DUMMY_3798 NETTRAN_DUMMY_3799 INV_X1 
XU1646 n529 n1521 NETTRAN_DUMMY_3800 NETTRAN_DUMMY_3801 INV_X1 
XU1645 n528 n1520 NETTRAN_DUMMY_3802 NETTRAN_DUMMY_3803 INV_X1 
XU1644 n551 n1501 NETTRAN_DUMMY_3804 NETTRAN_DUMMY_3805 INV_X1 
XU1643 n569 n1500 NETTRAN_DUMMY_3806 NETTRAN_DUMMY_3807 INV_X1 
XU1642 n535 n1499 NETTRAN_DUMMY_3808 NETTRAN_DUMMY_3809 INV_X1 
XU1641 n593 n1352 NETTRAN_DUMMY_3810 NETTRAN_DUMMY_3811 INV_X1 
XU1640 n524 n1333 NETTRAN_DUMMY_3812 NETTRAN_DUMMY_3813 INV_X1 
XU1639 n520 n1318 NETTRAN_DUMMY_3814 NETTRAN_DUMMY_3815 INV_X1 
XU1638 n515 n516 NETTRAN_DUMMY_3816 NETTRAN_DUMMY_3817 INV_X1 
XU1634 addr[0] n512 NETTRAN_DUMMY_3818 NETTRAN_DUMMY_3819 INV_X2 
XU1623 n500 n501 NETTRAN_DUMMY_3820 NETTRAN_DUMMY_3821 INV_X2 
XU1804 n12 n1536 NETTRAN_DUMMY_3822 NETTRAN_DUMMY_3823 INV_X1 
XU1803 n567 n1535 NETTRAN_DUMMY_3824 NETTRAN_DUMMY_3825 INV_X1 
XU1802 n565 n1534 NETTRAN_DUMMY_3826 NETTRAN_DUMMY_3827 INV_X1 
XU1801 n563 n1533 NETTRAN_DUMMY_3828 NETTRAN_DUMMY_3829 INV_X1 
XU1800 n612 n1532 NETTRAN_DUMMY_3830 NETTRAN_DUMMY_3831 INV_X1 
XU1799 n9 n1531 NETTRAN_DUMMY_3832 NETTRAN_DUMMY_3833 INV_X1 
XU1798 n629 n1530 NETTRAN_DUMMY_3834 NETTRAN_DUMMY_3835 INV_X1 
XU1797 n628 n1529 NETTRAN_DUMMY_3836 NETTRAN_DUMMY_3837 INV_X1 
XU1796 n531 n1528 NETTRAN_DUMMY_3838 NETTRAN_DUMMY_3839 INV_X1 
XU1795 n2 n1527 NETTRAN_DUMMY_3840 NETTRAN_DUMMY_3841 INV_X1 
XU1794 n45 n1851 NETTRAN_DUMMY_3842 NETTRAN_DUMMY_3843 INV_X1 
XU1793 n12 n493 n166 NETTRAN_DUMMY_3844 NETTRAN_DUMMY_3845 NAND2_X1 
XU1792 n1515 n1819 NETTRAN_DUMMY_3846 NETTRAN_DUMMY_3847 INV_X1 
XU1791 n413 n1651 NETTRAN_DUMMY_3848 NETTRAN_DUMMY_3849 INV_X1 
XU1790 n1506 n1801 NETTRAN_DUMMY_3850 NETTRAN_DUMMY_3851 INV_X1 
XU1789 n1160 n472 n1159 NETTRAN_DUMMY_3852 NETTRAN_DUMMY_3853 AND2_X1 
XU1788 n1084 n472 n1083 NETTRAN_DUMMY_3854 NETTRAN_DUMMY_3855 AND2_X1 
XU1787 n1825 n472 n1291 NETTRAN_DUMMY_3856 NETTRAN_DUMMY_3857 AND2_X1 
XU1786 n523 n444 n660 NETTRAN_DUMMY_3858 NETTRAN_DUMMY_3859 AND2_X1 
XU1785 n1501 n434 n1143 NETTRAN_DUMMY_3860 NETTRAN_DUMMY_3861 NAND2_X1 
XU1784 n513 n434 n431 NETTRAN_DUMMY_3862 NETTRAN_DUMMY_3863 AND2_X1 
XU1783 n1531 n449 n430 NETTRAN_DUMMY_3864 NETTRAN_DUMMY_3865 NOR2_X1 
XU1782 n1354 n472 n1353 NETTRAN_DUMMY_3866 NETTRAN_DUMMY_3867 AND2_X1 
XU1781 n1501 n461 n1190 NETTRAN_DUMMY_3868 NETTRAN_DUMMY_3869 NAND2_X1 
XU1780 n503 n1669 n1192 NETTRAN_DUMMY_3870 NETTRAN_DUMMY_3871 NOR2_X1 
XU1779 n1027 n472 n1026 NETTRAN_DUMMY_3872 NETTRAN_DUMMY_3873 AND2_X1 
XU1778 n884 n461 n883 NETTRAN_DUMMY_3874 NETTRAN_DUMMY_3875 AND2_X1 
XU1777 n765 n472 n764 NETTRAN_DUMMY_3876 NETTRAN_DUMMY_3877 AND2_X1 
XU1776 n565 n461 n566 n675 NETTRAN_DUMMY_3878 NETTRAN_DUMMY_3879 OAI21_X1 
XU1775 n1540 n493 n146 NETTRAN_DUMMY_3880 NETTRAN_DUMMY_3881 NOR2_X1 
XU1774 n551 n434 n1137 NETTRAN_DUMMY_3882 NETTRAN_DUMMY_3883 NAND2_X1 
XU1773 n431 n501 n433 n513 n1139 NETTRAN_DUMMY_3884 NETTRAN_DUMMY_3885 OAI22_X1 
XU1772 n536 n461 n1112 NETTRAN_DUMMY_3886 NETTRAN_DUMMY_3887 NOR2_X1 
XU1771 n574 n1665 NETTRAN_DUMMY_3888 NETTRAN_DUMMY_3889 INV_X1 
XU1770 n1545 n461 n689 NETTRAN_DUMMY_3890 NETTRAN_DUMMY_3891 NOR2_X1 
XU1769 n837 n444 n565 n836 NETTRAN_DUMMY_3892 NETTRAN_DUMMY_3893 OAI21_X1 
XU1768 n525 n461 n1668 n449 n759 NETTRAN_DUMMY_3894 NETTRAN_DUMMY_3895 OAI22_X1 
XU1767 n497 n439 n759 n758 NETTRAN_DUMMY_3896 NETTRAN_DUMMY_3897 AOI21_X1 
XU1766 n513 n445 n714 NETTRAN_DUMMY_3898 NETTRAN_DUMMY_3899 NOR2_X1 
XU1765 n1538 n497 n580 NETTRAN_DUMMY_3900 NETTRAN_DUMMY_3901 NOR2_X1 
XU1764 n461 n580 n1500 n501 n740 NETTRAN_DUMMY_3902 NETTRAN_DUMMY_3903 OAI22_X1 
XU1763 n855 n472 n854 NETTRAN_DUMMY_3904 NETTRAN_DUMMY_3905 AND2_X1 
XU1762 n551 n1849 n461 n1429 NETTRAN_DUMMY_3906 NETTRAN_DUMMY_3907 OAI21_X1 
XU1761 n1497 n1816 NETTRAN_DUMMY_3908 NETTRAN_DUMMY_3909 INV_X1 
XU1760 n488 n492 n429 NETTRAN_DUMMY_3910 NETTRAN_DUMMY_3911 XNOR2_X1 
XU1759 n548 n444 n597 NETTRAN_DUMMY_3912 NETTRAN_DUMMY_3913 NOR2_X1 
XU1758 n791 n792 n796 NETTRAN_DUMMY_3914 NETTRAN_DUMMY_3915 NOR2_X1 
XU1757 n1521 n434 n1133 NETTRAN_DUMMY_3916 NETTRAN_DUMMY_3917 NOR2_X1 
XU1756 n568 n664 n665 NETTRAN_DUMMY_3918 NETTRAN_DUMMY_3919 NOR2_X1 
XU1755 n461 n507 n428 NETTRAN_DUMMY_3920 NETTRAN_DUMMY_3921 XNOR2_X1 
XU1754 n1500 n472 n1498 NETTRAN_DUMMY_3922 NETTRAN_DUMMY_3923 NAND2_X1 
XU1753 n1687 n449 n448 n1682 n1707 NETTRAN_DUMMY_3924 NETTRAN_DUMMY_3925 AOI22_X1 
XU1752 n1707 n1688 N4640 NETTRAN_DUMMY_3926 NETTRAN_DUMMY_3927 NOR2_X1 
XU1751 n201 n444 n200 NETTRAN_DUMMY_3928 NETTRAN_DUMMY_3929 AND2_X1 
XU1750 n480 n449 n188 NETTRAN_DUMMY_3930 NETTRAN_DUMMY_3931 NOR2_X1 
XU1749 n434 n547 n546 NETTRAN_DUMMY_3932 NETTRAN_DUMMY_3933 NAND2_X1 
XU1748 n451 n1527 n16 NETTRAN_DUMMY_3934 NETTRAN_DUMMY_3935 NAND2_X1 
XU1747 n12 n1646 n488 n193 NETTRAN_DUMMY_3936 NETTRAN_DUMMY_3937 OAI21_X1 
XU1746 n539 n1778 n434 n994 NETTRAN_DUMMY_3938 NETTRAN_DUMMY_3939 OAI21_X1 
XU1745 n53 n437 n48 n259 NETTRAN_DUMMY_3940 NETTRAN_DUMMY_3941 OAI21_X1 
XU1744 n130 n437 n1643 n267 NETTRAN_DUMMY_3942 NETTRAN_DUMMY_3943 OAI21_X1 
XU1743 n817 n444 n1541 n816 NETTRAN_DUMMY_3944 NETTRAN_DUMMY_3945 OAI21_X1 
XU1742 n1771 n444 n1521 n807 NETTRAN_DUMMY_3946 NETTRAN_DUMMY_3947 OAI21_X1 
XU1741 n1774 n1534 n461 n1061 NETTRAN_DUMMY_3948 NETTRAN_DUMMY_3949 OAI21_X1 
XU1740 n36 n13 n488 n211 NETTRAN_DUMMY_3950 NETTRAN_DUMMY_3951 OAI21_X1 
XU1739 n593 n1501 n472 n873 NETTRAN_DUMMY_3952 NETTRAN_DUMMY_3953 OAI21_X1 
XU1738 n1783 n472 n1543 n967 NETTRAN_DUMMY_3954 NETTRAN_DUMMY_3955 OAI21_X1 
XU1737 n62 n1601 NETTRAN_DUMMY_3956 NETTRAN_DUMMY_3957 INV_X1 
XU1736 n130 n488 n1601 n129 NETTRAN_DUMMY_3958 NETTRAN_DUMMY_3959 OAI21_X1 
XU1735 n1499 n472 n1514 NETTRAN_DUMMY_3960 NETTRAN_DUMMY_3961 NAND2_X1 
XU1734 n1518 n1751 NETTRAN_DUMMY_3962 NETTRAN_DUMMY_3963 INV_X1 
XU1733 n1509 n1799 NETTRAN_DUMMY_3964 NETTRAN_DUMMY_3965 INV_X1 
XU1732 n1504 n1671 NETTRAN_DUMMY_3966 NETTRAN_DUMMY_3967 INV_X1 
XU1731 n1507 n1818 NETTRAN_DUMMY_3968 NETTRAN_DUMMY_3969 INV_X1 
XU1730 n6 n449 n427 NETTRAN_DUMMY_3970 NETTRAN_DUMMY_3971 AND2_X1 
XU1729 n493 n516 n604 NETTRAN_DUMMY_3972 NETTRAN_DUMMY_3973 NAND2_X1 
XU1728 n460 n21 n426 NETTRAN_DUMMY_3974 NETTRAN_DUMMY_3975 NAND2_X1 
XU1727 n1525 n516 n592 NETTRAN_DUMMY_3976 NETTRAN_DUMMY_3977 NAND2_X1 
XU1726 n1 n451 n407 NETTRAN_DUMMY_3978 NETTRAN_DUMMY_3979 NAND2_X1 
XU1725 n1531 n449 n406 NETTRAN_DUMMY_3980 NETTRAN_DUMMY_3981 NAND2_X1 
XU1724 n493 n1702 n1705 NETTRAN_DUMMY_3982 NETTRAN_DUMMY_3983 NOR2_X1 
XU1723 n434 n1664 n1705 n487 n1703 NETTRAN_DUMMY_3984 NETTRAN_DUMMY_3985 OAI211_X1 
XU1722 n1703 n1704 n1590 n434 N4680 NETTRAN_DUMMY_3986 NETTRAN_DUMMY_3987 OAI211_X1 
XU1721 n480 n461 n486 n1701 n1711 NETTRAN_DUMMY_3988 NETTRAN_DUMMY_3989 OAI22_X1 
XU1720 n1712 n497 n1709 NETTRAN_DUMMY_3990 NETTRAN_DUMMY_3991 OR2_X1 
XU1719 n1699 n497 n1711 n512 n1710 NETTRAN_DUMMY_3992 NETTRAN_DUMMY_3993 NAND4_X1 
XU1718 n433 n1709 n1710 N19750 NETTRAN_DUMMY_3994 NETTRAN_DUMMY_3995 AOI21_X1 
XU1717 n449 n1540 n11 NETTRAN_DUMMY_3996 NETTRAN_DUMMY_3997 NAND2_X1 
XU1716 n1537 n449 n55 NETTRAN_DUMMY_3998 NETTRAN_DUMMY_3999 NAND2_X1 
XU1715 n29 n484 n11 n306 NETTRAN_DUMMY_4000 NETTRAN_DUMMY_4001 AOI21_X1 
XU1714 n18 n484 n36 n205 NETTRAN_DUMMY_4002 NETTRAN_DUMMY_4003 AOI21_X1 
XU1713 n488 n204 n203 NETTRAN_DUMMY_4004 NETTRAN_DUMMY_4005 NAND2_X1 
XU1712 IN0 n487 n1727 n1728 n1718 NETTRAN_DUMMY_4006 NETTRAN_DUMMY_4007 OAI211_X1 
XU1849 n445 n472 n520 n712 NETTRAN_DUMMY_4008 NETTRAN_DUMMY_4009 AND3_X1 
XU1823 n434 n1682 n1699 n1524 N19520 NETTRAN_DUMMY_4010 NETTRAN_DUMMY_4011 AND4_X1 
XU1822 n444 n488 n38 n207 NETTRAN_DUMMY_4012 NETTRAN_DUMMY_4013 NAND3_X1 
XU1821 n449 n512 n52 NETTRAN_DUMMY_4014 NETTRAN_DUMMY_4015 NAND2_X1 
XU1820 n512 n1682 n1713 NETTRAN_DUMMY_4016 NETTRAN_DUMMY_4017 NAND2_X1 
XU1819 n445 n493 n823 NETTRAN_DUMMY_4018 NETTRAN_DUMMY_4019 NOR2_X1 
XU1818 n484 n449 n14 NETTRAN_DUMMY_4020 NETTRAN_DUMMY_4021 NAND2_X1 
XU1817 n497 n472 n624 NETTRAN_DUMMY_4022 NETTRAN_DUMMY_4023 NAND2_X1 
XU1816 n480 n493 n1524 n1737 NETTRAN_DUMMY_4024 NETTRAN_DUMMY_4025 NAND3_X1 
XU1815 n1737 n480 n1708 n1735 NETTRAN_DUMMY_4026 NETTRAN_DUMMY_4027 OAI21_X1 
XU1814 n1684 n1524 n472 n1733 NETTRAN_DUMMY_4028 NETTRAN_DUMMY_4029 AOI21_X1 
XU1813 n513 n488 n434 n1722 NETTRAN_DUMMY_4030 NETTRAN_DUMMY_4031 AOI21_X1 
XU1812 n497 n461 n480 n1724 NETTRAN_DUMMY_4032 NETTRAN_DUMMY_4033 NAND3_X1 
XU1811 n445 n434 n1704 NETTRAN_DUMMY_4034 NETTRAN_DUMMY_4035 NAND2_X1 
XU1810 n1524 n493 n1740 NETTRAN_DUMMY_4036 NETTRAN_DUMMY_4037 NAND2_X1 
XU1809 n433 n497 IN0 n480 n1740 n1738 NETTRAN_DUMMY_4038 NETTRAN_DUMMY_4039 AOI221_X1 
XU1808 n1589 n1586 n1739 NETTRAN_DUMMY_4040 NETTRAN_DUMMY_4041 NOR2_X1 
XU1807 n1739 n463 n1738 n452 n461 N13181 NETTRAN_DUMMY_4042 NETTRAN_DUMMY_4043 OAI221_X1 
XU1806 n501 n449 n12 NETTRAN_DUMMY_4044 NETTRAN_DUMMY_4045 NAND2_X1 
XU1805 n1684 n461 n434 n1727 NETTRAN_DUMMY_4046 NETTRAN_DUMMY_4047 NOR3_X1 
XCLKBUF_X1_G2B1I1 clk n63_G2B1I1 NETTRAN_DUMMY_4048 NETTRAN_DUMMY_4049 CLKBUF_X1 
XCLKBUF_X1_G2B1I3 clk n63_G2B1I3 NETTRAN_DUMMY_4050 NETTRAN_DUMMY_4051 CLKBUF_X1 
XCLKBUF_X1_G2B1I4 clk n63_G2B1I4 NETTRAN_DUMMY_4052 NETTRAN_DUMMY_4053 CLKBUF_X1 
XCLKBUF_X1_G2B1I5 clk n63_G2B1I5 NETTRAN_DUMMY_4054 NETTRAN_DUMMY_4055 CLKBUF_X1 
XCLKBUF_X1_G2B1I7 clk n63_G2B1I7 NETTRAN_DUMMY_4056 NETTRAN_DUMMY_4057 CLKBUF_X1 
XCLKBUF_X1_G2B1I9 clk n63_G2B1I9 NETTRAN_DUMMY_4058 NETTRAN_DUMMY_4059 CLKBUF_X1 
XCLKBUF_X1_G2B1I6 clk n63_G2B1I6 NETTRAN_DUMMY_4060 NETTRAN_DUMMY_4061 CLKBUF_X1 
XU14 n468 n463 NETTRAN_DUMMY_4062 NETTRAN_DUMMY_4063 BUF_X1 
XU47 d[29] n457 NETTRAN_DUMMY_4064 NETTRAN_DUMMY_4065 BUF_X1 
XU483 N19750 n459 NETTRAN_DUMMY_4066 NETTRAN_DUMMY_4067 BUF_X16 
XU485 d[9] n465 NETTRAN_DUMMY_4068 NETTRAN_DUMMY_4069 INV_X1 
XU494 n465 n467 NETTRAN_DUMMY_4070 NETTRAN_DUMMY_4071 INV_X32 
XU498 d[8] n469 NETTRAN_DUMMY_4072 NETTRAN_DUMMY_4073 INV_X1 
XU513 n469 n470 NETTRAN_DUMMY_4074 NETTRAN_DUMMY_4075 INV_X16 
XU532 d[6] n474 NETTRAN_DUMMY_4076 NETTRAN_DUMMY_4077 BUF_X1 
XU585 d[5] n476 NETTRAN_DUMMY_4078 NETTRAN_DUMMY_4079 INV_X1 
XU773 n476 n478 NETTRAN_DUMMY_4080 NETTRAN_DUMMY_4081 INV_X16 
XU1590 n1856 n479 NETTRAN_DUMMY_4082 NETTRAN_DUMMY_4083 INV_X1 
XU1592 n479 n481 NETTRAN_DUMMY_4084 NETTRAN_DUMMY_4085 INV_X8 
XU1593 N4870 n482 NETTRAN_DUMMY_4086 NETTRAN_DUMMY_4087 INV_X1 
XU1594 n482 n483 NETTRAN_DUMMY_4088 NETTRAN_DUMMY_4089 INV_X8 
XU1596 n468 n485 NETTRAN_DUMMY_4090 NETTRAN_DUMMY_4091 INV_X1 
XU1599 n485 n486 NETTRAN_DUMMY_4092 NETTRAN_DUMMY_4093 INV_X16 
XU1604 N5090 n489 NETTRAN_DUMMY_4094 NETTRAN_DUMMY_4095 INV_X1 
XU1618 n489 n490 NETTRAN_DUMMY_4096 NETTRAN_DUMMY_4097 INV_X32 
XU1620 d[48] n491 NETTRAN_DUMMY_4098 NETTRAN_DUMMY_4099 INV_X1 
XU1626 n491 n494 NETTRAN_DUMMY_4100 NETTRAN_DUMMY_4101 INV_X32 
XU1627 d[47] n496 NETTRAN_DUMMY_4102 NETTRAN_DUMMY_4103 BUF_X1 
XU1628 d[46] n498 NETTRAN_DUMMY_4104 NETTRAN_DUMMY_4105 BUF_X1 
XU1630 d[45] n504 NETTRAN_DUMMY_4106 NETTRAN_DUMMY_4107 BUF_X1 
XU1632 d[44] n505 NETTRAN_DUMMY_4108 NETTRAN_DUMMY_4109 INV_X1 
XU1633 n505 n506 NETTRAN_DUMMY_4110 NETTRAN_DUMMY_4111 INV_X16 
XU1636 N13181 n508 NETTRAN_DUMMY_4112 NETTRAN_DUMMY_4113 INV_X1 
XU1833 n508 n510 NETTRAN_DUMMY_4114 NETTRAN_DUMMY_4115 INV_X32 
XU1835 N13331 n511 NETTRAN_DUMMY_4116 NETTRAN_DUMMY_4117 INV_X1 
XU1836 n511 n514 NETTRAN_DUMMY_4118 NETTRAN_DUMMY_4119 INV_X32 
XU1837 N13521 n1546 NETTRAN_DUMMY_4120 NETTRAN_DUMMY_4121 INV_X32 
XU1838 n1546 n1548 NETTRAN_DUMMY_4122 NETTRAN_DUMMY_4123 INV_X1 
XU1839 n2010 n1549 NETTRAN_DUMMY_4124 NETTRAN_DUMMY_4125 CLKBUF_X1 
XU1840 n1551 n1550 NETTRAN_DUMMY_4126 NETTRAN_DUMMY_4127 CLKBUF_X1 
XU1841 n1549 n1551 NETTRAN_DUMMY_4128 NETTRAN_DUMMY_4129 INV_X32 
XU1842 n1550 c2[16] NETTRAN_DUMMY_4130 NETTRAN_DUMMY_4131 INV_X32 
XU1843 n2009 n1553 NETTRAN_DUMMY_4132 NETTRAN_DUMMY_4133 CLKBUF_X1 
XU1844 n1555 n1554 NETTRAN_DUMMY_4134 NETTRAN_DUMMY_4135 CLKBUF_X1 
XU1845 n1553 n1555 NETTRAN_DUMMY_4136 NETTRAN_DUMMY_4137 INV_X32 
XU1846 n1554 c2[15] NETTRAN_DUMMY_4138 NETTRAN_DUMMY_4139 INV_X32 
XU1847 n2008 n1557 NETTRAN_DUMMY_4140 NETTRAN_DUMMY_4141 CLKBUF_X1 
XU1848 n1559 n1558 NETTRAN_DUMMY_4142 NETTRAN_DUMMY_4143 CLKBUF_X1 
XU1850 n1557 n1559 NETTRAN_DUMMY_4144 NETTRAN_DUMMY_4145 INV_X32 
XU1851 n1558 c2[14] NETTRAN_DUMMY_4146 NETTRAN_DUMMY_4147 INV_X32 
XU1852 n2007 n1561 NETTRAN_DUMMY_4148 NETTRAN_DUMMY_4149 CLKBUF_X1 
XU1853 n1563 n1562 NETTRAN_DUMMY_4150 NETTRAN_DUMMY_4151 CLKBUF_X1 
XU1854 n1561 n1563 NETTRAN_DUMMY_4152 NETTRAN_DUMMY_4153 INV_X32 
XU1855 n1562 c2[13] NETTRAN_DUMMY_4154 NETTRAN_DUMMY_4155 INV_X32 
XU1856 n2006 n1565 NETTRAN_DUMMY_4156 NETTRAN_DUMMY_4157 CLKBUF_X1 
XU1857 n1567 n1566 NETTRAN_DUMMY_4158 NETTRAN_DUMMY_4159 CLKBUF_X1 
XU1858 n1565 n1567 NETTRAN_DUMMY_4160 NETTRAN_DUMMY_4161 INV_X32 
XU1859 n1566 c2[12] NETTRAN_DUMMY_4162 NETTRAN_DUMMY_4163 INV_X32 
XU1860 n2018 n1569 NETTRAN_DUMMY_4164 NETTRAN_DUMMY_4165 CLKBUF_X1 
XU1861 n1571 n1570 NETTRAN_DUMMY_4166 NETTRAN_DUMMY_4167 CLKBUF_X1 
XU1862 n1569 n1571 NETTRAN_DUMMY_4168 NETTRAN_DUMMY_4169 INV_X32 
XU1863 n1570 c2[11] NETTRAN_DUMMY_4170 NETTRAN_DUMMY_4171 INV_X32 
XU1864 n2017 n1573 NETTRAN_DUMMY_4172 NETTRAN_DUMMY_4173 CLKBUF_X1 
XU1865 n1575 n1574 NETTRAN_DUMMY_4174 NETTRAN_DUMMY_4175 CLKBUF_X1 
XU1866 n1573 n1575 NETTRAN_DUMMY_4176 NETTRAN_DUMMY_4177 INV_X32 
XU1867 n1574 c2[10] NETTRAN_DUMMY_4178 NETTRAN_DUMMY_4179 INV_X32 
XU1868 n2016 n1577 NETTRAN_DUMMY_4180 NETTRAN_DUMMY_4181 CLKBUF_X1 
XU1869 n1579 n1578 NETTRAN_DUMMY_4182 NETTRAN_DUMMY_4183 CLKBUF_X1 
XU1870 n1577 n1579 NETTRAN_DUMMY_4184 NETTRAN_DUMMY_4185 INV_X32 
XU1871 n1578 c2[9] NETTRAN_DUMMY_4186 NETTRAN_DUMMY_4187 INV_X32 
XU1872 n2015 n1581 NETTRAN_DUMMY_4188 NETTRAN_DUMMY_4189 CLKBUF_X1 
XU1873 n1583 n1582 NETTRAN_DUMMY_4190 NETTRAN_DUMMY_4191 CLKBUF_X1 
XU1874 n1581 n1583 NETTRAN_DUMMY_4192 NETTRAN_DUMMY_4193 INV_X32 
XU1875 n1582 c2[8] NETTRAN_DUMMY_4194 NETTRAN_DUMMY_4195 INV_X32 
XU1876 n2014 n1592 NETTRAN_DUMMY_4196 NETTRAN_DUMMY_4197 CLKBUF_X1 
XU1877 n1764 n1750 NETTRAN_DUMMY_4198 NETTRAN_DUMMY_4199 CLKBUF_X1 
XU1878 n1592 n1764 NETTRAN_DUMMY_4200 NETTRAN_DUMMY_4201 INV_X32 
XU1879 n1750 c2[7] NETTRAN_DUMMY_4202 NETTRAN_DUMMY_4203 INV_X32 
XU1880 n2013 n1782 NETTRAN_DUMMY_4204 NETTRAN_DUMMY_4205 CLKBUF_X1 
XU1881 n1788 n1786 NETTRAN_DUMMY_4206 NETTRAN_DUMMY_4207 CLKBUF_X1 
XU1882 n1782 n1788 NETTRAN_DUMMY_4208 NETTRAN_DUMMY_4209 INV_X32 
XU1883 n1786 c2[6] NETTRAN_DUMMY_4210 NETTRAN_DUMMY_4211 INV_X32 
XU1884 n2012 n1793 NETTRAN_DUMMY_4212 NETTRAN_DUMMY_4213 CLKBUF_X1 
XU1885 n1798 n1794 NETTRAN_DUMMY_4214 NETTRAN_DUMMY_4215 CLKBUF_X1 
XU1886 n1793 n1798 NETTRAN_DUMMY_4216 NETTRAN_DUMMY_4217 INV_X32 
XU1887 n1794 c2[5] NETTRAN_DUMMY_4218 NETTRAN_DUMMY_4219 INV_X32 
XU1888 n2011 n1802 NETTRAN_DUMMY_4220 NETTRAN_DUMMY_4221 CLKBUF_X1 
XU1889 n1807 n1803 NETTRAN_DUMMY_4222 NETTRAN_DUMMY_4223 CLKBUF_X1 
XU1890 n1802 n1807 NETTRAN_DUMMY_4224 NETTRAN_DUMMY_4225 INV_X32 
XU1891 n1803 c2[4] NETTRAN_DUMMY_4226 NETTRAN_DUMMY_4227 INV_X32 
XU1892 n2026 n1810 NETTRAN_DUMMY_4228 NETTRAN_DUMMY_4229 CLKBUF_X1 
XU1893 n1820 n1813 NETTRAN_DUMMY_4230 NETTRAN_DUMMY_4231 CLKBUF_X1 
XU1894 n1810 n1820 NETTRAN_DUMMY_4232 NETTRAN_DUMMY_4233 INV_X32 
XU1895 n1813 c2[3] NETTRAN_DUMMY_4234 NETTRAN_DUMMY_4235 INV_X32 
XU1896 n2025 n1823 NETTRAN_DUMMY_4236 NETTRAN_DUMMY_4237 CLKBUF_X1 
XU1897 n1830 n1829 NETTRAN_DUMMY_4238 NETTRAN_DUMMY_4239 CLKBUF_X1 
XU1898 n1823 n1830 NETTRAN_DUMMY_4240 NETTRAN_DUMMY_4241 INV_X32 
XU1899 n1829 c2[2] NETTRAN_DUMMY_4242 NETTRAN_DUMMY_4243 INV_X32 
XU1900 n2024 n1837 NETTRAN_DUMMY_4244 NETTRAN_DUMMY_4245 CLKBUF_X1 
XU1901 n1854 n1843 NETTRAN_DUMMY_4246 NETTRAN_DUMMY_4247 CLKBUF_X1 
XU1902 n1837 n1854 NETTRAN_DUMMY_4248 NETTRAN_DUMMY_4249 INV_X32 
XU1903 n1843 c2[1] NETTRAN_DUMMY_4250 NETTRAN_DUMMY_4251 INV_X32 
XU1904 n2023 n1858 NETTRAN_DUMMY_4252 NETTRAN_DUMMY_4253 CLKBUF_X1 
XU1905 n1860 n1859 NETTRAN_DUMMY_4254 NETTRAN_DUMMY_4255 CLKBUF_X1 
XU1906 n1858 n1860 NETTRAN_DUMMY_4256 NETTRAN_DUMMY_4257 INV_X32 
XU1907 n1859 c2[0] NETTRAN_DUMMY_4258 NETTRAN_DUMMY_4259 INV_X32 
XU1908 n2058 n1862 NETTRAN_DUMMY_4260 NETTRAN_DUMMY_4261 CLKBUF_X1 
XU1909 n1864 n1863 NETTRAN_DUMMY_4262 NETTRAN_DUMMY_4263 CLKBUF_X1 
XU1910 n1862 n1864 NETTRAN_DUMMY_4264 NETTRAN_DUMMY_4265 INV_X32 
XU1911 n1863 c0[7] NETTRAN_DUMMY_4266 NETTRAN_DUMMY_4267 INV_X32 
XU1912 n2057 n1866 NETTRAN_DUMMY_4268 NETTRAN_DUMMY_4269 CLKBUF_X1 
XU1913 n1868 n1867 NETTRAN_DUMMY_4270 NETTRAN_DUMMY_4271 CLKBUF_X1 
XU1914 n1866 n1868 NETTRAN_DUMMY_4272 NETTRAN_DUMMY_4273 INV_X32 
XU1915 n1867 c0[6] NETTRAN_DUMMY_4274 NETTRAN_DUMMY_4275 INV_X32 
XU1916 n2056 n1870 NETTRAN_DUMMY_4276 NETTRAN_DUMMY_4277 CLKBUF_X1 
XU1917 n1872 n1871 NETTRAN_DUMMY_4278 NETTRAN_DUMMY_4279 CLKBUF_X1 
XU1918 n1870 n1872 NETTRAN_DUMMY_4280 NETTRAN_DUMMY_4281 INV_X32 
XU1919 n1871 c0[5] NETTRAN_DUMMY_4282 NETTRAN_DUMMY_4283 INV_X32 
XU1920 n2055 n1874 NETTRAN_DUMMY_4284 NETTRAN_DUMMY_4285 CLKBUF_X1 
XU1921 n1876 n1875 NETTRAN_DUMMY_4286 NETTRAN_DUMMY_4287 CLKBUF_X1 
XU1922 n1874 n1876 NETTRAN_DUMMY_4288 NETTRAN_DUMMY_4289 INV_X32 
XU1923 n1875 c0[4] NETTRAN_DUMMY_4290 NETTRAN_DUMMY_4291 INV_X32 
XU1924 n2054 n1878 NETTRAN_DUMMY_4292 NETTRAN_DUMMY_4293 CLKBUF_X1 
XU1925 n1880 n1879 NETTRAN_DUMMY_4294 NETTRAN_DUMMY_4295 CLKBUF_X1 
XU1926 n1878 n1880 NETTRAN_DUMMY_4296 NETTRAN_DUMMY_4297 INV_X32 
XU1927 n1879 c0[3] NETTRAN_DUMMY_4298 NETTRAN_DUMMY_4299 INV_X32 
XU1928 n2053 n1882 NETTRAN_DUMMY_4300 NETTRAN_DUMMY_4301 CLKBUF_X1 
XU1929 n1884 n1883 NETTRAN_DUMMY_4302 NETTRAN_DUMMY_4303 CLKBUF_X1 
XU1930 n1882 n1884 NETTRAN_DUMMY_4304 NETTRAN_DUMMY_4305 INV_X32 
XU1931 n1883 c0[2] NETTRAN_DUMMY_4306 NETTRAN_DUMMY_4307 INV_X32 
XU1932 n2052 n1886 NETTRAN_DUMMY_4308 NETTRAN_DUMMY_4309 CLKBUF_X1 
XU1933 n1888 n1887 NETTRAN_DUMMY_4310 NETTRAN_DUMMY_4311 CLKBUF_X1 
XU1934 n1886 n1888 NETTRAN_DUMMY_4312 NETTRAN_DUMMY_4313 INV_X32 
XU1935 n1887 c0[1] NETTRAN_DUMMY_4314 NETTRAN_DUMMY_4315 INV_X32 
XU1936 n2051 n1890 NETTRAN_DUMMY_4316 NETTRAN_DUMMY_4317 CLKBUF_X1 
XU1937 n1892 n1891 NETTRAN_DUMMY_4318 NETTRAN_DUMMY_4319 CLKBUF_X1 
XU1938 n1890 n1892 NETTRAN_DUMMY_4320 NETTRAN_DUMMY_4321 INV_X32 
XU1939 n1891 c0[0] NETTRAN_DUMMY_4322 NETTRAN_DUMMY_4323 INV_X32 
XU1940 n2022 n1894 NETTRAN_DUMMY_4324 NETTRAN_DUMMY_4325 CLKBUF_X1 
XU1941 n1896 n1895 NETTRAN_DUMMY_4326 NETTRAN_DUMMY_4327 CLKBUF_X1 
XU1942 n1894 n1896 NETTRAN_DUMMY_4328 NETTRAN_DUMMY_4329 INV_X32 
XU1943 n1895 c1[17] NETTRAN_DUMMY_4330 NETTRAN_DUMMY_4331 INV_X32 
XU1944 n2021 n1898 NETTRAN_DUMMY_4332 NETTRAN_DUMMY_4333 CLKBUF_X1 
XU1945 n1900 n1899 NETTRAN_DUMMY_4334 NETTRAN_DUMMY_4335 CLKBUF_X1 
XU1946 n1898 n1900 NETTRAN_DUMMY_4336 NETTRAN_DUMMY_4337 INV_X32 
XU1947 n1899 c1[16] NETTRAN_DUMMY_4338 NETTRAN_DUMMY_4339 INV_X32 
XU1948 n2020 n1902 NETTRAN_DUMMY_4340 NETTRAN_DUMMY_4341 CLKBUF_X1 
XU1949 n1904 n1903 NETTRAN_DUMMY_4342 NETTRAN_DUMMY_4343 CLKBUF_X1 
XU1950 n1902 n1904 NETTRAN_DUMMY_4344 NETTRAN_DUMMY_4345 INV_X32 
XU1951 n1903 c1[15] NETTRAN_DUMMY_4346 NETTRAN_DUMMY_4347 INV_X32 
XU1952 n2019 n1906 NETTRAN_DUMMY_4348 NETTRAN_DUMMY_4349 CLKBUF_X1 
XU1953 n1908 n1907 NETTRAN_DUMMY_4350 NETTRAN_DUMMY_4351 CLKBUF_X1 
XU1954 n1906 n1908 NETTRAN_DUMMY_4352 NETTRAN_DUMMY_4353 INV_X32 
XU1955 n1907 c1[14] NETTRAN_DUMMY_4354 NETTRAN_DUMMY_4355 INV_X32 
XU1956 n2034 n1910 NETTRAN_DUMMY_4356 NETTRAN_DUMMY_4357 CLKBUF_X1 
XU1957 n1912 n1911 NETTRAN_DUMMY_4358 NETTRAN_DUMMY_4359 CLKBUF_X1 
XU1958 n1910 n1912 NETTRAN_DUMMY_4360 NETTRAN_DUMMY_4361 INV_X32 
XU1959 n1911 c1[13] NETTRAN_DUMMY_4362 NETTRAN_DUMMY_4363 INV_X32 
XU1960 n2033 n1914 NETTRAN_DUMMY_4364 NETTRAN_DUMMY_4365 CLKBUF_X1 
XU1961 n1916 n1915 NETTRAN_DUMMY_4366 NETTRAN_DUMMY_4367 CLKBUF_X1 
XU1962 n1914 n1916 NETTRAN_DUMMY_4368 NETTRAN_DUMMY_4369 INV_X32 
XU1963 n1915 c1[12] NETTRAN_DUMMY_4370 NETTRAN_DUMMY_4371 INV_X32 
XU1964 n1921 c1[11] NETTRAN_DUMMY_4372 NETTRAN_DUMMY_4373 BUF_X1 
XU1965 n1920 n1919 NETTRAN_DUMMY_4374 NETTRAN_DUMMY_4375 CLKBUF_X1 
XU1966 n2032 n1920 NETTRAN_DUMMY_4376 NETTRAN_DUMMY_4377 INV_X32 
XU1967 n1919 n1921 NETTRAN_DUMMY_4378 NETTRAN_DUMMY_4379 INV_X32 
XU1968 n2031 n1922 NETTRAN_DUMMY_4380 NETTRAN_DUMMY_4381 CLKBUF_X1 
XU1969 n1924 n1923 NETTRAN_DUMMY_4382 NETTRAN_DUMMY_4383 CLKBUF_X1 
XU1970 n1922 n1924 NETTRAN_DUMMY_4384 NETTRAN_DUMMY_4385 INV_X32 
XU1971 n1923 c1[10] NETTRAN_DUMMY_4386 NETTRAN_DUMMY_4387 INV_X32 
XU1972 n2030 n1926 NETTRAN_DUMMY_4388 NETTRAN_DUMMY_4389 CLKBUF_X1 
XU1973 n1928 n1927 NETTRAN_DUMMY_4390 NETTRAN_DUMMY_4391 CLKBUF_X1 
XU1974 n1926 n1928 NETTRAN_DUMMY_4392 NETTRAN_DUMMY_4393 INV_X32 
XU1975 n1927 c1[9] NETTRAN_DUMMY_4394 NETTRAN_DUMMY_4395 INV_X32 
XU1976 n2029 n1930 NETTRAN_DUMMY_4396 NETTRAN_DUMMY_4397 CLKBUF_X1 
XU1977 n1932 n1931 NETTRAN_DUMMY_4398 NETTRAN_DUMMY_4399 CLKBUF_X1 
XU1978 n1930 n1932 NETTRAN_DUMMY_4400 NETTRAN_DUMMY_4401 INV_X32 
XU1979 n1931 c1[8] NETTRAN_DUMMY_4402 NETTRAN_DUMMY_4403 INV_X32 
XU1980 n1937 c1[7] NETTRAN_DUMMY_4404 NETTRAN_DUMMY_4405 BUF_X1 
XU1981 n1936 n1935 NETTRAN_DUMMY_4406 NETTRAN_DUMMY_4407 CLKBUF_X1 
XU1982 n2028 n1936 NETTRAN_DUMMY_4408 NETTRAN_DUMMY_4409 INV_X32 
XU1983 n1935 n1937 NETTRAN_DUMMY_4410 NETTRAN_DUMMY_4411 INV_X32 
XU1984 n2027 n1938 NETTRAN_DUMMY_4412 NETTRAN_DUMMY_4413 CLKBUF_X1 
XU1985 n1940 n1939 NETTRAN_DUMMY_4414 NETTRAN_DUMMY_4415 CLKBUF_X1 
XU1986 n1938 n1940 NETTRAN_DUMMY_4416 NETTRAN_DUMMY_4417 INV_X32 
XU1987 n1939 c1[6] NETTRAN_DUMMY_4418 NETTRAN_DUMMY_4419 INV_X32 
XU1988 n2042 n1942 NETTRAN_DUMMY_4420 NETTRAN_DUMMY_4421 CLKBUF_X1 
XU1989 n1944 n1943 NETTRAN_DUMMY_4422 NETTRAN_DUMMY_4423 CLKBUF_X1 
XU1990 n1942 n1944 NETTRAN_DUMMY_4424 NETTRAN_DUMMY_4425 INV_X32 
XU1991 n1943 c1[5] NETTRAN_DUMMY_4426 NETTRAN_DUMMY_4427 INV_X32 
XU1992 n2041 n1946 NETTRAN_DUMMY_4428 NETTRAN_DUMMY_4429 CLKBUF_X1 
XU1993 n1948 n1947 NETTRAN_DUMMY_4430 NETTRAN_DUMMY_4431 CLKBUF_X1 
XU1994 n1946 n1948 NETTRAN_DUMMY_4432 NETTRAN_DUMMY_4433 INV_X32 
XU1995 n1947 c1[4] NETTRAN_DUMMY_4434 NETTRAN_DUMMY_4435 INV_X32 
XU1996 n2040 n1950 NETTRAN_DUMMY_4436 NETTRAN_DUMMY_4437 CLKBUF_X1 
XU1997 n1952 n1951 NETTRAN_DUMMY_4438 NETTRAN_DUMMY_4439 CLKBUF_X1 
XU1998 n1950 n1952 NETTRAN_DUMMY_4440 NETTRAN_DUMMY_4441 INV_X32 
XU1999 n1951 c1[3] NETTRAN_DUMMY_4442 NETTRAN_DUMMY_4443 INV_X32 
XU2000 n1957 c1[2] NETTRAN_DUMMY_4444 NETTRAN_DUMMY_4445 BUF_X1 
XU2001 n1956 n1955 NETTRAN_DUMMY_4446 NETTRAN_DUMMY_4447 CLKBUF_X1 
XU2002 n2039 n1956 NETTRAN_DUMMY_4448 NETTRAN_DUMMY_4449 INV_X32 
XU2003 n1955 n1957 NETTRAN_DUMMY_4450 NETTRAN_DUMMY_4451 INV_X32 
XU2004 n2038 n1958 NETTRAN_DUMMY_4452 NETTRAN_DUMMY_4453 CLKBUF_X1 
XU2005 n1960 n1959 NETTRAN_DUMMY_4454 NETTRAN_DUMMY_4455 CLKBUF_X1 
XU2006 n1958 n1960 NETTRAN_DUMMY_4456 NETTRAN_DUMMY_4457 INV_X32 
XU2007 n1959 c1[1] NETTRAN_DUMMY_4458 NETTRAN_DUMMY_4459 INV_X32 
XU2008 n2037 n1962 NETTRAN_DUMMY_4460 NETTRAN_DUMMY_4461 CLKBUF_X1 
XU2009 n1964 n1963 NETTRAN_DUMMY_4462 NETTRAN_DUMMY_4463 CLKBUF_X1 
XU2010 n1962 n1964 NETTRAN_DUMMY_4464 NETTRAN_DUMMY_4465 INV_X32 
XU2011 n1963 c1[0] NETTRAN_DUMMY_4466 NETTRAN_DUMMY_4467 INV_X32 
XU2012 n2036 n1966 NETTRAN_DUMMY_4468 NETTRAN_DUMMY_4469 CLKBUF_X1 
XU2013 n1968 n1967 NETTRAN_DUMMY_4470 NETTRAN_DUMMY_4471 CLKBUF_X1 
XU2014 n1966 n1968 NETTRAN_DUMMY_4472 NETTRAN_DUMMY_4473 INV_X32 
XU2015 n1967 c0[17] NETTRAN_DUMMY_4474 NETTRAN_DUMMY_4475 INV_X32 
XU2016 n2035 n1970 NETTRAN_DUMMY_4476 NETTRAN_DUMMY_4477 CLKBUF_X1 
XU2017 n1972 n1971 NETTRAN_DUMMY_4478 NETTRAN_DUMMY_4479 CLKBUF_X1 
XU2018 n1970 n1972 NETTRAN_DUMMY_4480 NETTRAN_DUMMY_4481 INV_X32 
XU2019 n1971 c0[16] NETTRAN_DUMMY_4482 NETTRAN_DUMMY_4483 INV_X32 
XU2020 n2050 n1974 NETTRAN_DUMMY_4484 NETTRAN_DUMMY_4485 CLKBUF_X1 
XU2021 n1976 n1975 NETTRAN_DUMMY_4486 NETTRAN_DUMMY_4487 CLKBUF_X1 
XU2022 n1974 n1976 NETTRAN_DUMMY_4488 NETTRAN_DUMMY_4489 INV_X32 
XU2023 n1975 c0[15] NETTRAN_DUMMY_4490 NETTRAN_DUMMY_4491 INV_X32 
XU2024 n2049 n1978 NETTRAN_DUMMY_4492 NETTRAN_DUMMY_4493 CLKBUF_X1 
XU2025 n1980 n1979 NETTRAN_DUMMY_4494 NETTRAN_DUMMY_4495 CLKBUF_X1 
XU2026 n1978 n1980 NETTRAN_DUMMY_4496 NETTRAN_DUMMY_4497 INV_X32 
XU2027 n1979 c0[14] NETTRAN_DUMMY_4498 NETTRAN_DUMMY_4499 INV_X32 
XU2028 n2048 n1982 NETTRAN_DUMMY_4500 NETTRAN_DUMMY_4501 CLKBUF_X1 
XU2029 n1984 n1983 NETTRAN_DUMMY_4502 NETTRAN_DUMMY_4503 CLKBUF_X1 
XU2030 n1982 n1984 NETTRAN_DUMMY_4504 NETTRAN_DUMMY_4505 INV_X32 
XU2031 n1983 c0[13] NETTRAN_DUMMY_4506 NETTRAN_DUMMY_4507 INV_X32 
XU2032 n1989 c0[12] NETTRAN_DUMMY_4508 NETTRAN_DUMMY_4509 BUF_X1 
XU2033 n1988 n1987 NETTRAN_DUMMY_4510 NETTRAN_DUMMY_4511 CLKBUF_X1 
XU2034 n2047 n1988 NETTRAN_DUMMY_4512 NETTRAN_DUMMY_4513 INV_X32 
XU2035 n1987 n1989 NETTRAN_DUMMY_4514 NETTRAN_DUMMY_4515 INV_X32 
XU2036 n2046 n1990 NETTRAN_DUMMY_4516 NETTRAN_DUMMY_4517 CLKBUF_X1 
XU2037 n1992 n1991 NETTRAN_DUMMY_4518 NETTRAN_DUMMY_4519 CLKBUF_X1 
XU2038 n1990 n1992 NETTRAN_DUMMY_4520 NETTRAN_DUMMY_4521 INV_X32 
XU2039 n1991 c0[11] NETTRAN_DUMMY_4522 NETTRAN_DUMMY_4523 INV_X32 
XU2040 n2045 n1994 NETTRAN_DUMMY_4524 NETTRAN_DUMMY_4525 CLKBUF_X1 
XU2041 n1996 n1995 NETTRAN_DUMMY_4526 NETTRAN_DUMMY_4527 CLKBUF_X1 
XU2042 n1994 n1996 NETTRAN_DUMMY_4528 NETTRAN_DUMMY_4529 INV_X32 
XU2043 n1995 c0[10] NETTRAN_DUMMY_4530 NETTRAN_DUMMY_4531 INV_X32 
XU2044 n2001 c0[9] NETTRAN_DUMMY_4532 NETTRAN_DUMMY_4533 BUF_X1 
XU2045 n2000 n1999 NETTRAN_DUMMY_4534 NETTRAN_DUMMY_4535 CLKBUF_X1 
XU2046 n2044 n2000 NETTRAN_DUMMY_4536 NETTRAN_DUMMY_4537 INV_X32 
XU2047 n1999 n2001 NETTRAN_DUMMY_4538 NETTRAN_DUMMY_4539 INV_X32 
XU2048 n2043 n2002 NETTRAN_DUMMY_4540 NETTRAN_DUMMY_4541 CLKBUF_X1 
XU2049 n2004 n2003 NETTRAN_DUMMY_4542 NETTRAN_DUMMY_4543 CLKBUF_X1 
XU2050 n2002 n2004 NETTRAN_DUMMY_4544 NETTRAN_DUMMY_4545 INV_X32 
XU2051 n2003 c0[8] NETTRAN_DUMMY_4546 NETTRAN_DUMMY_4547 INV_X32 
XU2052 n409 n2059 NETTRAN_DUMMY_4548 NETTRAN_DUMMY_4549 BUF_X1 
XU2053 n483 n2060 NETTRAN_DUMMY_4550 NETTRAN_DUMMY_4551 BUF_X1 
XU2054 n510 n2061 NETTRAN_DUMMY_4552 NETTRAN_DUMMY_4553 BUF_X1 
.ENDS

.SUBCKT gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff clk rstn ce valid_out 
+ IN0 IN1 data_out[63] data_out[62] data_out[61] data_out[60] data_out[59] data_out[58] 
+ data_out[57] data_out[56] data_out[55] data_out[54] data_out[53] data_out[52] 
+ data_out[51] data_out[50] data_out[49] data_out[48] data_out[47] data_out[46] 
+ data_out[45] data_out[44] data_out[43] data_out[42] data_out[41] data_out[40] 
+ data_out[39] data_out[38] data_out[37] data_out[36] data_out[35] data_out[34] 
+ data_out[33] data_out[32] data_out[31] data_out[30] data_out[29] data_out[28] 
+ data_out[27] data_out[26] data_out[25] data_out[24] data_out[23] data_out[22] 
+ data_out[21] data_out[20] data_out[19] data_out[18] data_out[17] data_out[16] 
+ data_out[15] data_out[14] data_out[13] data_out[12] data_out[11] data_out[10] 
+ data_out[9] data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] data_out[3] 
+ data_out[2] data_out[1] data_out[0] IN2 IN3 clk_cts_3 
Xz1_reg_3_ n748 n84_G2B1I5 z1_next[27] n121 NETTRAN_DUMMY_4554 NETTRAN_DUMMY_4555 DFF_X1 
Xz1_reg_42_ n2007 n78_G2B1I8 z1[42] n79 NETTRAN_DUMMY_4556 NETTRAN_DUMMY_4557 DFF_X1 
Xz1_reg_18_ n1997 n84 z1_next[42] n106 NETTRAN_DUMMY_4558 NETTRAN_DUMMY_4559 DFF_X1 
Xz1_reg_52_ n747 n78_G2B1I8 z1[52] n67 NETTRAN_DUMMY_4560 NETTRAN_DUMMY_4561 DFF_X1 
Xz1_reg_28_ n746 n84_G2B1I3 z1_next[52] n96 NETTRAN_DUMMY_4562 NETTRAN_DUMMY_4563 DFF_X1 
Xz1_reg_4_ n745 n76_G2B1I4 z1_next[28] n120 NETTRAN_DUMMY_4564 NETTRAN_DUMMY_4565 DFF_X1 
Xz1_reg_43_ n1976 n84_G2B1I4 z1[43] n77 NETTRAN_DUMMY_4566 NETTRAN_DUMMY_4567 DFF_X1 
Xz1_reg_19_ n744 n84_G2B1I3 z1_next[43] n105 NETTRAN_DUMMY_4568 NETTRAN_DUMMY_4569 DFF_X1 
Xz1_reg_53_ n742 n84_G2B1I3 z1[53] n66 NETTRAN_DUMMY_4570 NETTRAN_DUMMY_4571 DFF_X1 
Xz1_reg_29_ n741 n76_G2B1I4 z1_next[53] n95 NETTRAN_DUMMY_4572 NETTRAN_DUMMY_4573 DFF_X1 
Xz1_reg_5_ n740 n76_G2B1I4 z1_next[29] n119 NETTRAN_DUMMY_4574 NETTRAN_DUMMY_4575 DFF_X1 
Xz1_reg_63_ n1949 n84_G2B1I3 NETTRAN_DUMMY_4576 n56 NETTRAN_DUMMY_4577 NETTRAN_DUMMY_4578 DFF_X1 
Xz1_reg_39_ n739 n84_G2B1I3 z1_next[63] n85 NETTRAN_DUMMY_4579 NETTRAN_DUMMY_4580 DFF_X1 
Xz1_reg_15_ n738 n84_G2B1I6 z1_next[39] n109 NETTRAN_DUMMY_4581 NETTRAN_DUMMY_4582 DFF_X1 
Xz1_reg_49_ n1933 n84_G2B1I6 z1[49] n70 NETTRAN_DUMMY_4583 NETTRAN_DUMMY_4584 DFF_X1 
Xz1_reg_25_ n734 n84_G2B1I4 z1_next[49] n99 NETTRAN_DUMMY_4585 NETTRAN_DUMMY_4586 DFF_X1 
Xz1_reg_1_ n1926 n84_G2B1I5 z1_next[25] n123 NETTRAN_DUMMY_4587 NETTRAN_DUMMY_4588 DFF_X1 
Xz3_reg_61_ n733 n82_G2B1I3 z3[61] n3 NETTRAN_DUMMY_4589 NETTRAN_DUMMY_4590 DFF_X1 
Xz3_reg_54_ n731 n82_G2B1I7 z3_next[61] n10 NETTRAN_DUMMY_4591 NETTRAN_DUMMY_4592 DFF_X1 
Xz3_reg_47_ n730 n82_G2B1I3 NETTRAN_DUMMY_4593 n17 NETTRAN_DUMMY_4594 NETTRAN_DUMMY_4595 DFF_X1 
Xz3_reg_40_ n728 n80_G2B1I6 NETTRAN_DUMMY_4596 n24 NETTRAN_DUMMY_4597 NETTRAN_DUMMY_4598 DFF_X1 
Xz3_reg_33_ n556 n80_G2B1I2 z3_next[40] n31 NETTRAN_DUMMY_4599 NETTRAN_DUMMY_4600 DFF_X1 
Xz3_reg_26_ n1896 n80_G2B1I6 z3_next[33] n38 NETTRAN_DUMMY_4601 NETTRAN_DUMMY_4602 DFF_X1 
Xz3_reg_19_ n1891 n80_G2B1I6 NETTRAN_DUMMY_4603 n45 NETTRAN_DUMMY_4604 NETTRAN_DUMMY_4605 DFF_X1 
Xz3_reg_12_ n724 n80_G2B1I2 z3_next[19] n52 NETTRAN_DUMMY_4606 NETTRAN_DUMMY_4607 DFF_X1 
Xz3_reg_57_ n1879 n82_G2B1I3 z3[57] n7 NETTRAN_DUMMY_4608 NETTRAN_DUMMY_4609 DFF_X1 
Xz3_reg_50_ n722 n82_G2B1I5 NETTRAN_DUMMY_4610 n14 NETTRAN_DUMMY_4611 NETTRAN_DUMMY_4612 DFF_X1 
Xz3_reg_43_ n721 n80_G2B1I2 NETTRAN_DUMMY_4613 n21 NETTRAN_DUMMY_4614 NETTRAN_DUMMY_4615 DFF_X1 
Xz3_reg_36_ n1861 n76_G2B1I1 z3_next[43] n28 NETTRAN_DUMMY_4616 NETTRAN_DUMMY_4617 DFF_X1 
Xz3_reg_29_ n720 n76_G2B1I4 z3_next[36] n35 NETTRAN_DUMMY_4618 NETTRAN_DUMMY_4619 DFF_X1 
Xz3_reg_22_ n718 n76_G2B1I3 NETTRAN_DUMMY_4620 n42 NETTRAN_DUMMY_4621 NETTRAN_DUMMY_4622 DFF_X1 
Xz3_reg_15_ n1849 n76_G2B1I3 z3_next[22] n49 NETTRAN_DUMMY_4623 NETTRAN_DUMMY_4624 DFF_X1 
Xz3_reg_60_ n717 n82_G2B1I4 z3[60] n4 NETTRAN_DUMMY_4625 NETTRAN_DUMMY_4626 DFF_X1 
Xz3_reg_53_ n1835 n84_G2B1I5 NETTRAN_DUMMY_4627 n11 NETTRAN_DUMMY_4628 NETTRAN_DUMMY_4629 DFF_X1 
Xz3_reg_46_ n716 n84_G2B1I5 NETTRAN_DUMMY_4630 n18 NETTRAN_DUMMY_4631 NETTRAN_DUMMY_4632 DFF_X1 
Xz3_reg_39_ n715 n84_G2B1I5 z3_next[46] n25 NETTRAN_DUMMY_4633 NETTRAN_DUMMY_4634 DFF_X1 
Xz3_reg_32_ n714 n84_G2B1I5 z3_next[39] n32 NETTRAN_DUMMY_4635 NETTRAN_DUMMY_4636 DFF_X1 
Xz3_reg_25_ n713 n80_G2B1I5 z3_next[32] n39 NETTRAN_DUMMY_4637 NETTRAN_DUMMY_4638 DFF_X1 
Xz3_reg_18_ n712 n84_G2B1I5 NETTRAN_DUMMY_4639 n46 NETTRAN_DUMMY_4640 NETTRAN_DUMMY_4641 DFF_X1 
Xz3_reg_11_ n1804 n84_G2B1I2 z3_next[18] n53 NETTRAN_DUMMY_4642 NETTRAN_DUMMY_4643 DFF_X1 
Xz3_reg_63_ n711 n84_G2B1I4 z3[63] n1 NETTRAN_DUMMY_4644 NETTRAN_DUMMY_4645 DFF_X1 
Xz3_reg_56_ n710 n82_G2B1I4 z3_next[63] n8 NETTRAN_DUMMY_4646 NETTRAN_DUMMY_4647 DFF_X1 
Xz3_reg_49_ n1787 clk_G1B1I2 NETTRAN_DUMMY_4648 n15 NETTRAN_DUMMY_4649 NETTRAN_DUMMY_4650 DFF_X1 
Xz3_reg_42_ n709 n82_G2B1I8 NETTRAN_DUMMY_4651 n22 NETTRAN_DUMMY_4652 NETTRAN_DUMMY_4653 DFF_X1 
Xz3_reg_35_ n708 n82_G2B1I7 z3_next[42] n29 NETTRAN_DUMMY_4654 NETTRAN_DUMMY_4655 DFF_X1 
Xz3_reg_28_ n1772 n82_G2B1I7 z3_next[35] n36 NETTRAN_DUMMY_4656 NETTRAN_DUMMY_4657 DFF_X1 
Xz3_reg_21_ n707 n82_G2B1I6 NETTRAN_DUMMY_4658 n43 NETTRAN_DUMMY_4659 NETTRAN_DUMMY_4660 DFF_X1 
Xz3_reg_14_ n705 n80_G2B1I6 z3_next[21] n50 NETTRAN_DUMMY_4661 NETTRAN_DUMMY_4662 DFF_X1 
Xz3_reg_59_ n704 n82_G2B1I3 z3[59] n5 NETTRAN_DUMMY_4663 NETTRAN_DUMMY_4664 DFF_X1 
Xz3_reg_52_ n702 n82_G2B1I3 NETTRAN_DUMMY_4665 n12 NETTRAN_DUMMY_4666 NETTRAN_DUMMY_4667 DFF_X1 
Xz3_reg_45_ n1750 n82_G2B1I6 NETTRAN_DUMMY_4668 n19 NETTRAN_DUMMY_4669 NETTRAN_DUMMY_4670 DFF_X1 
Xz3_reg_38_ n1745 n82_G2B1I6 z3_next[45] n26 NETTRAN_DUMMY_4671 NETTRAN_DUMMY_4672 DFF_X1 
Xz3_reg_31_ n1740 n82_G2B1I5 z3_next[38] n33 NETTRAN_DUMMY_4673 NETTRAN_DUMMY_4674 DFF_X1 
Xz3_reg_24_ n1731 n76_G2B1I1 z3_next[31] n40 NETTRAN_DUMMY_4675 NETTRAN_DUMMY_4676 DFF_X1 
Xz3_reg_17_ n697 n76_G2B1I1 z3_next[24] n47 NETTRAN_DUMMY_4677 NETTRAN_DUMMY_4678 DFF_X1 
Xz3_reg_10_ n1724 n76_G2B1I1 z3_next[17] n54 NETTRAN_DUMMY_4679 NETTRAN_DUMMY_4680 DFF_X1 
Xz3_reg_62_ n1717 n82_G2B1I3 z3[62] n2 NETTRAN_DUMMY_4681 NETTRAN_DUMMY_4682 DFF_X1 
Xz3_reg_55_ n695 n82_G2B1I7 z3_next[62] n9 NETTRAN_DUMMY_4683 NETTRAN_DUMMY_4684 DFF_X1 
Xz3_reg_48_ n1704 n82_G2B1I7 NETTRAN_DUMMY_4685 n16 NETTRAN_DUMMY_4686 NETTRAN_DUMMY_4687 DFF_X1 
Xz3_reg_41_ n694 n82_G2B1I7 NETTRAN_DUMMY_4688 n23 NETTRAN_DUMMY_4689 NETTRAN_DUMMY_4690 DFF_X1 
Xz3_reg_34_ n693 n82_G2B1I7 z3_next[41] n30 NETTRAN_DUMMY_4691 NETTRAN_DUMMY_4692 DFF_X1 
Xz3_reg_27_ n1688 n82_G2B1I5 z3_next[34] n37 NETTRAN_DUMMY_4693 NETTRAN_DUMMY_4694 DFF_X1 
Xz3_reg_20_ n692 n82_G2B1I6 NETTRAN_DUMMY_4695 n44 NETTRAN_DUMMY_4696 NETTRAN_DUMMY_4697 DFF_X1 
Xz3_reg_13_ n690 n80_G2B1I6 z3_next[20] n51 NETTRAN_DUMMY_4698 NETTRAN_DUMMY_4699 DFF_X1 
Xz3_reg_58_ n688 n82_G2B1I7 z3[58] n6 NETTRAN_DUMMY_4700 NETTRAN_DUMMY_4701 DFF_X1 
Xz3_reg_51_ n687 n82_G2B1I5 z3_next[58] n13 NETTRAN_DUMMY_4702 NETTRAN_DUMMY_4703 DFF_X1 
Xz3_reg_44_ n686 n82_G2B1I6 NETTRAN_DUMMY_4704 n20 NETTRAN_DUMMY_4705 NETTRAN_DUMMY_4706 DFF_X1 
Xz3_reg_37_ n685 n82_G2B1I6 z3_next[44] n27 NETTRAN_DUMMY_4707 NETTRAN_DUMMY_4708 DFF_X1 
Xz3_reg_30_ n684 n82_G2B1I8 z3_next[37] n34 NETTRAN_DUMMY_4709 NETTRAN_DUMMY_4710 DFF_X1 
Xz3_reg_23_ n683 n76_G2B1I3 NETTRAN_DUMMY_4711 n41 NETTRAN_DUMMY_4712 NETTRAN_DUMMY_4713 DFF_X1 
Xz3_reg_16_ n1644 n76 z3_next[23] n48 NETTRAN_DUMMY_4714 NETTRAN_DUMMY_4715 DFF_X1 
Xz3_reg_9_ n681 n76_G2B1I1 z3_next[16] n55 NETTRAN_DUMMY_4716 NETTRAN_DUMMY_4717 DFF_X1 
XU22 n188 n261 NETTRAN_DUMMY_4718 NETTRAN_DUMMY_4719 BUF_X2 
XU21 n188 n260 NETTRAN_DUMMY_4720 NETTRAN_DUMMY_4721 BUF_X2 
XU20 n188 n259 NETTRAN_DUMMY_4722 NETTRAN_DUMMY_4723 BUF_X2 
XU16 n255 n256 NETTRAN_DUMMY_4724 NETTRAN_DUMMY_4725 INV_X1 
XU12 rstn n252 NETTRAN_DUMMY_4726 NETTRAN_DUMMY_4727 INV_X1 
XU11 IN0 n250 NETTRAN_DUMMY_4728 NETTRAN_DUMMY_4729 INV_X1 
XU10 IN1 n248 NETTRAN_DUMMY_4730 NETTRAN_DUMMY_4731 INV_X1 
XU9 IN3 n246 NETTRAN_DUMMY_4732 NETTRAN_DUMMY_4733 INV_X1 
XU7 IN2 n185 NETTRAN_DUMMY_4734 NETTRAN_DUMMY_4735 INV_X1 
Xz2_reg_24_ n1631 n82_G2B1I4 z2_next[37] n166 NETTRAN_DUMMY_4736 NETTRAN_DUMMY_4737 DFF_X1 
Xz2_reg_11_ n1625 n82_G2B1I4 z2_next[24] n179 NETTRAN_DUMMY_4738 NETTRAN_DUMMY_4739 DFF_X1 
Xz2_reg_56_ n680 n76_G2B1I1 NETTRAN_DUMMY_4740 n134 NETTRAN_DUMMY_4741 NETTRAN_DUMMY_4742 DFF_X1 
Xz2_reg_43_ n679 n76_G2B1I1 z2_next[56] n147 NETTRAN_DUMMY_4743 NETTRAN_DUMMY_4744 DFF_X1 
Xz2_reg_30_ n678 n76_G2B1I1 z2_next[43] n160 NETTRAN_DUMMY_4745 NETTRAN_DUMMY_4746 DFF_X1 
Xz2_reg_17_ n1604 n76_G2B1I3 z2_next[30] n173 NETTRAN_DUMMY_4747 NETTRAN_DUMMY_4748 DFF_X1 
Xz2_reg_62_ n677 n125_G2B1I3 z2[62] n126 NETTRAN_DUMMY_4749 NETTRAN_DUMMY_4750 DFF_X1 
Xz2_reg_49_ n675 n82_G2B1I8 z2_next[62] n141 NETTRAN_DUMMY_4751 NETTRAN_DUMMY_4752 DFF_X1 
Xz2_reg_36_ n674 n125_G2B1I3 z2_next[49] n154 NETTRAN_DUMMY_4753 NETTRAN_DUMMY_4754 DFF_X1 
Xz2_reg_23_ n1587 n76_G2B1I3 z2_next[36] n167 NETTRAN_DUMMY_4755 NETTRAN_DUMMY_4756 DFF_X1 
Xz2_reg_10_ n1577 n76 z2_next[23] n180 NETTRAN_DUMMY_4757 NETTRAN_DUMMY_4758 DFF_X1 
Xz2_reg_55_ n672 n125_G2B1I3 NETTRAN_DUMMY_4759 n135 NETTRAN_DUMMY_4760 NETTRAN_DUMMY_4761 DFF_X1 
Xz2_reg_42_ n1565 n76 z2_next[55] n148 NETTRAN_DUMMY_4762 NETTRAN_DUMMY_4763 DFF_X1 
Xz2_reg_29_ n1560 n76_G2B1I4 z2_next[42] n161 NETTRAN_DUMMY_4764 NETTRAN_DUMMY_4765 DFF_X1 
Xz2_reg_16_ n1554 n76_G2B1I3 z2_next[29] n174 NETTRAN_DUMMY_4766 NETTRAN_DUMMY_4767 DFF_X1 
Xz2_reg_61_ n671 n125_G2B1I3 z2[61] n128 NETTRAN_DUMMY_4768 NETTRAN_DUMMY_4769 DFF_X1 
Xz2_reg_48_ n669 n82_G2B1I8 z2_next[61] n142 NETTRAN_DUMMY_4770 NETTRAN_DUMMY_4771 DFF_X1 
Xz2_reg_35_ n668 n82_G2B1I8 z2_next[48] n155 NETTRAN_DUMMY_4772 NETTRAN_DUMMY_4773 DFF_X1 
Xz2_reg_22_ n1535 clk_G1B1I2 z2_next[35] n168 NETTRAN_DUMMY_4774 NETTRAN_DUMMY_4775 DFF_X1 
Xz2_reg_9_ n666 n76_G2B1I1 z2_next[22] n181 NETTRAN_DUMMY_4776 NETTRAN_DUMMY_4777 DFF_X1 
Xz2_reg_54_ n665 n82_G2B1I8 NETTRAN_DUMMY_4778 n136 NETTRAN_DUMMY_4779 NETTRAN_DUMMY_4780 DFF_X1 
Xz2_reg_41_ n663 clk_G1B1I2 z2_next[54] n149 NETTRAN_DUMMY_4781 NETTRAN_DUMMY_4782 DFF_X1 
Xz2_reg_28_ n662 n82_G2B1I5 z2_next[41] n162 NETTRAN_DUMMY_4783 NETTRAN_DUMMY_4784 DFF_X1 
Xz2_reg_15_ n661 n82_G2B1I5 z2_next[28] n175 NETTRAN_DUMMY_4785 NETTRAN_DUMMY_4786 DFF_X1 
Xz2_reg_60_ n659 n82_G2B1I5 NETTRAN_DUMMY_4787 n130 NETTRAN_DUMMY_4788 NETTRAN_DUMMY_4789 DFF_X1 
Xz2_reg_47_ n658 n80_G2B1I2 z2_next[60] n143 NETTRAN_DUMMY_4790 NETTRAN_DUMMY_4791 DFF_X1 
Xz2_reg_34_ n657 n80_G2B1I7 z2_next[47] n156 NETTRAN_DUMMY_4792 NETTRAN_DUMMY_4793 DFF_X1 
Xz2_reg_21_ n656 n80_G2B1I7 z2_next[34] n169 NETTRAN_DUMMY_4794 NETTRAN_DUMMY_4795 DFF_X1 
Xz2_reg_8_ n1482 n80_G2B1I7 z2_next[21] n182 NETTRAN_DUMMY_4796 NETTRAN_DUMMY_4797 DFF_X1 
Xz2_reg_53_ n654 n80_G2B1I4 NETTRAN_DUMMY_4798 n137 NETTRAN_DUMMY_4799 NETTRAN_DUMMY_4800 DFF_X1 
Xz2_reg_40_ n653 n80_G2B1I5 z2_next[53] n150 NETTRAN_DUMMY_4801 NETTRAN_DUMMY_4802 DFF_X1 
Xz2_reg_27_ n651 n80_G2B1I5 z2_next[40] n163 NETTRAN_DUMMY_4803 NETTRAN_DUMMY_4804 DFF_X1 
Xz2_reg_14_ n1461 n80_G2B1I6 z2_next[27] n176 NETTRAN_DUMMY_4805 NETTRAN_DUMMY_4806 DFF_X1 
Xz2_reg_59_ n650 n80_G2B1I4 NETTRAN_DUMMY_4807 n131 NETTRAN_DUMMY_4808 NETTRAN_DUMMY_4809 DFF_X1 
Xz2_reg_46_ n1450 n80_G2B1I6 z2_next[59] n144 NETTRAN_DUMMY_4810 NETTRAN_DUMMY_4811 DFF_X1 
Xz2_reg_33_ n649 n80_G2B1I1 z2_next[46] n157 NETTRAN_DUMMY_4812 NETTRAN_DUMMY_4813 DFF_X1 
Xz2_reg_20_ n1439 n80_G2B1I7 z2_next[33] n170 NETTRAN_DUMMY_4814 NETTRAN_DUMMY_4815 DFF_X1 
Xz2_reg_7_ n648 n80_G2B1I1 z2_next[20] n183 NETTRAN_DUMMY_4816 NETTRAN_DUMMY_4817 DFF_X1 
Xz2_reg_52_ n647 n80_G2B1I4 NETTRAN_DUMMY_4818 n138 NETTRAN_DUMMY_4819 NETTRAN_DUMMY_4820 DFF_X1 
Xz2_reg_39_ n646 n80_G2B1I2 z2_next[52] n151 NETTRAN_DUMMY_4821 NETTRAN_DUMMY_4822 DFF_X1 
Xz2_reg_26_ n1422 n80 z2_next[39] n164 NETTRAN_DUMMY_4823 NETTRAN_DUMMY_4824 DFF_X1 
Xz2_reg_13_ n1412 n80 z2_next[26] n177 NETTRAN_DUMMY_4825 NETTRAN_DUMMY_4826 DFF_X1 
Xz2_reg_58_ n645 n80_G2B1I4 NETTRAN_DUMMY_4827 n132 NETTRAN_DUMMY_4828 NETTRAN_DUMMY_4829 DFF_X1 
Xz2_reg_45_ n642 n80_G2B1I1 z2_next[58] n145 NETTRAN_DUMMY_4830 NETTRAN_DUMMY_4831 DFF_X1 
Xz2_reg_32_ n1401 n80_G2B1I7 z2_next[45] n158 NETTRAN_DUMMY_4832 NETTRAN_DUMMY_4833 DFF_X1 
Xz2_reg_19_ n641 n80_G2B1I1 z2_next[32] n171 NETTRAN_DUMMY_4834 NETTRAN_DUMMY_4835 DFF_X1 
Xz2_reg_6_ n1387 n80_G2B1I5 z2_next[19] n184 NETTRAN_DUMMY_4836 NETTRAN_DUMMY_4837 DFF_X1 
Xz1_reg_59_ n639 n78_G2B1I7 NETTRAN_DUMMY_4838 n60 NETTRAN_DUMMY_4839 NETTRAN_DUMMY_4840 DFF_X1 
Xz1_reg_35_ n638 n80_G2B1I1 z1_next[59] n89 NETTRAN_DUMMY_4841 NETTRAN_DUMMY_4842 DFF_X1 
Xz1_reg_11_ n636 n78_G2B1I6 z1_next[35] n113 NETTRAN_DUMMY_4843 NETTRAN_DUMMY_4844 DFF_X1 
Xz1_reg_45_ n635 n78_G2B1I6 z1[45] n74 NETTRAN_DUMMY_4845 NETTRAN_DUMMY_4846 DFF_X1 
Xz1_reg_21_ n634 n78_G2B1I6 z1_next[45] n103 NETTRAN_DUMMY_4847 NETTRAN_DUMMY_4848 DFF_X1 
Xz1_reg_60_ n633 n78_G2B1I6 NETTRAN_DUMMY_4849 n59 NETTRAN_DUMMY_4850 NETTRAN_DUMMY_4851 DFF_X1 
Xz1_reg_36_ n632 n78_G2B1I7 z1_next[60] n88 NETTRAN_DUMMY_4852 NETTRAN_DUMMY_4853 DFF_X1 
Xz1_reg_12_ n630 n78_G2B1I4 z1_next[36] n112 NETTRAN_DUMMY_4854 NETTRAN_DUMMY_4855 DFF_X1 
Xz1_reg_55_ n629 n78_G2B1I2 NETTRAN_DUMMY_4856 n64 NETTRAN_DUMMY_4857 NETTRAN_DUMMY_4858 DFF_X1 
Xz1_reg_31_ n628 n84_G2B1I6 z1_next[55] n93 NETTRAN_DUMMY_4859 NETTRAN_DUMMY_4860 DFF_X1 
Xz1_reg_7_ n627 n84_G2B1I6 z1_next[31] n117 NETTRAN_DUMMY_4861 NETTRAN_DUMMY_4862 DFF_X1 
Xz1_reg_46_ n617 n78_G2B1I4 z1[46] n73 NETTRAN_DUMMY_4863 NETTRAN_DUMMY_4864 DFF_X1 
Xz1_reg_22_ n616 n78_G2B1I5 z1_next[46] n102 NETTRAN_DUMMY_4865 NETTRAN_DUMMY_4866 DFF_X1 
Xz1_reg_61_ n615 n78_G2B1I5 NETTRAN_DUMMY_4867 n58 NETTRAN_DUMMY_4868 NETTRAN_DUMMY_4869 DFF_X1 
Xz1_reg_37_ n614 n78_G2B1I2 z1_next[61] n87 NETTRAN_DUMMY_4870 NETTRAN_DUMMY_4871 DFF_X1 
Xz1_reg_13_ n613 n78_G2B1I4 z1_next[37] n111 NETTRAN_DUMMY_4872 NETTRAN_DUMMY_4873 DFF_X1 
Xz1_reg_56_ n611 n78_G2B1I8 NETTRAN_DUMMY_4874 n63 NETTRAN_DUMMY_4875 NETTRAN_DUMMY_4876 DFF_X1 
Xz1_reg_32_ n608 n78_G2B1I8 z1_next[56] n92 NETTRAN_DUMMY_4877 NETTRAN_DUMMY_4878 DFF_X1 
Xz1_reg_8_ n1295 n78_G2B1I8 z1_next[32] n116 NETTRAN_DUMMY_4879 NETTRAN_DUMMY_4880 DFF_X1 
Xz1_reg_47_ n607 n78_G2B1I8 z1[47] n72 NETTRAN_DUMMY_4881 NETTRAN_DUMMY_4882 DFF_X1 
Xz1_reg_23_ n606 n78_G2B1I5 z1_next[47] n101 NETTRAN_DUMMY_4883 NETTRAN_DUMMY_4884 DFF_X1 
Xz1_reg_62_ n605 n84 NETTRAN_DUMMY_4885 n57 NETTRAN_DUMMY_4886 NETTRAN_DUMMY_4887 DFF_X1 
Xz1_reg_38_ n604 n84_G2B1I4 z1_next[62] n86 NETTRAN_DUMMY_4888 NETTRAN_DUMMY_4889 DFF_X1 
Xz1_reg_14_ n602 n84_G2B1I6 z1_next[38] n110 NETTRAN_DUMMY_4890 NETTRAN_DUMMY_4891 DFF_X1 
Xz1_reg_57_ n1261 n78_G2B1I8 NETTRAN_DUMMY_4892 n62 NETTRAN_DUMMY_4893 NETTRAN_DUMMY_4894 DFF_X1 
Xz1_reg_33_ n601 n78_G2B1I2 z1_next[57] n91 NETTRAN_DUMMY_4895 NETTRAN_DUMMY_4896 DFF_X1 
Xz1_reg_9_ n1250 n78_G2B1I2 z1_next[33] n115 NETTRAN_DUMMY_4897 NETTRAN_DUMMY_4898 DFF_X1 
Xz1_reg_48_ n599 n84_G2B1I4 z1[48] n71 NETTRAN_DUMMY_4899 NETTRAN_DUMMY_4900 DFF_X1 
Xz1_reg_24_ n598 n76_G2B1I4 z1_next[48] n100 NETTRAN_DUMMY_4901 NETTRAN_DUMMY_4902 DFF_X1 
Xz1_reg_58_ n1234 n84 NETTRAN_DUMMY_4903 n61 NETTRAN_DUMMY_4904 NETTRAN_DUMMY_4905 DFF_X1 
Xz1_reg_34_ n596 n78_G2B1I2 NETTRAN_DUMMY_4906 n90 NETTRAN_DUMMY_4907 NETTRAN_DUMMY_4908 DFF_X1 
Xz1_reg_10_ n1228 n78_G2B1I7 z1_next[34] n114 NETTRAN_DUMMY_4909 NETTRAN_DUMMY_4910 DFF_X1 
Xz1_reg_44_ n594 n84_G2B1I6 z1[44] n75 NETTRAN_DUMMY_4911 NETTRAN_DUMMY_4912 DFF_X1 
Xz1_reg_20_ n593 n84_G2B1I6 z1_next[44] n104 NETTRAN_DUMMY_4913 NETTRAN_DUMMY_4914 DFF_X1 
Xz1_reg_54_ n591 n84 z1[54] n65 NETTRAN_DUMMY_4915 NETTRAN_DUMMY_4916 DFF_X1 
Xz1_reg_30_ n590 n84_G2B1I3 z1_next[54] n94 NETTRAN_DUMMY_4917 NETTRAN_DUMMY_4918 DFF_X1 
Xz1_reg_6_ n589 n84_G2B1I3 z1_next[30] n118 NETTRAN_DUMMY_4919 NETTRAN_DUMMY_4920 DFF_X1 
Xz1_reg_40_ n588 n80_G2B1I7 z1[40] n83 NETTRAN_DUMMY_4921 NETTRAN_DUMMY_4922 DFF_X1 
Xz1_reg_16_ n586 n78_G2B1I6 z1_next[40] n108 NETTRAN_DUMMY_4923 NETTRAN_DUMMY_4924 DFF_X1 
Xz1_reg_50_ n584 n78_G2B1I7 z1[50] n69 NETTRAN_DUMMY_4925 NETTRAN_DUMMY_4926 DFF_X1 
Xz1_reg_26_ n583 n80_G2B1I5 z1_next[50] n98 NETTRAN_DUMMY_4927 NETTRAN_DUMMY_4928 DFF_X1 
Xz1_reg_2_ n582 n80_G2B1I5 z1_next[26] n122 NETTRAN_DUMMY_4929 NETTRAN_DUMMY_4930 DFF_X1 
Xz1_reg_41_ n1169 n78_G2B1I7 z1[41] n81 NETTRAN_DUMMY_4931 NETTRAN_DUMMY_4932 DFF_X1 
Xz1_reg_17_ n581 n78_G2B1I6 z1_next[41] n107 NETTRAN_DUMMY_4933 NETTRAN_DUMMY_4934 DFF_X1 
Xz1_reg_51_ n578 n78_G2B1I4 z1[51] n68 NETTRAN_DUMMY_4935 NETTRAN_DUMMY_4936 DFF_X1 
Xz1_reg_27_ n577 n84_G2B1I6 z1_next[51] n97 NETTRAN_DUMMY_4937 NETTRAN_DUMMY_4938 DFF_X1 
XU422 n197 n216 n340 NETTRAN_DUMMY_4939 NETTRAN_DUMMY_4940 XOR2_X1 
XU421 n231 n340 n339 NETTRAN_DUMMY_4941 NETTRAN_DUMMY_4942 XOR2_X1 
XU420 n74 z1[50] n215 NETTRAN_DUMMY_4943 NETTRAN_DUMMY_4944 XOR2_X1 
XU419 n196 n215 n338 NETTRAN_DUMMY_4945 NETTRAN_DUMMY_4946 XOR2_X1 
XU418 n230 n338 n337 NETTRAN_DUMMY_4947 NETTRAN_DUMMY_4948 XOR2_X1 
XU417 n73 z1[51] n214 NETTRAN_DUMMY_4949 NETTRAN_DUMMY_4950 XOR2_X1 
XU416 n195 n214 n336 NETTRAN_DUMMY_4951 NETTRAN_DUMMY_4952 XOR2_X1 
XU415 n229 n336 n335 NETTRAN_DUMMY_4953 NETTRAN_DUMMY_4954 XOR2_X1 
XU414 n72 z1[52] n213 NETTRAN_DUMMY_4955 NETTRAN_DUMMY_4956 XOR2_X1 
XU413 n194 n213 n334 NETTRAN_DUMMY_4957 NETTRAN_DUMMY_4958 XOR2_X1 
XU412 n228 n334 n333 NETTRAN_DUMMY_4959 NETTRAN_DUMMY_4960 XOR2_X1 
XU411 n71 z1[53] n212 NETTRAN_DUMMY_4961 NETTRAN_DUMMY_4962 XOR2_X1 
XU410 n193 n212 n332 NETTRAN_DUMMY_4963 NETTRAN_DUMMY_4964 XOR2_X1 
XU409 n227 n332 n331 NETTRAN_DUMMY_4965 NETTRAN_DUMMY_4966 XOR2_X1 
XU408 n70 z1[54] n211 NETTRAN_DUMMY_4967 NETTRAN_DUMMY_4968 XOR2_X1 
XU407 n192 n211 n330 NETTRAN_DUMMY_4969 NETTRAN_DUMMY_4970 XOR2_X1 
XU406 n226 n330 n329 NETTRAN_DUMMY_4971 NETTRAN_DUMMY_4972 XOR2_X1 
Xdata_out_reg_0_ n555 n125_G2B1I6 n2025 NETTRAN_DUMMY_4973 NETTRAN_DUMMY_4974 NETTRAN_DUMMY_4975 DFF_X1 
Xdata_out_reg_1_ n1142 n78_G2B1I5 data_out[1] NETTRAN_DUMMY_4976 NETTRAN_DUMMY_4977 
+ NETTRAN_DUMMY_4978 DFF_X1 
Xdata_out_reg_2_ n1137 n82_G2B1I3 data_out[2] NETTRAN_DUMMY_4979 NETTRAN_DUMMY_4980 
+ NETTRAN_DUMMY_4981 DFF_X1 
Xdata_out_reg_3_ n1132 n82_G2B1I2 data_out[3] NETTRAN_DUMMY_4982 NETTRAN_DUMMY_4983 
+ NETTRAN_DUMMY_4984 DFF_X1 
Xdata_out_reg_4_ n1127 n82_G2B1I2 data_out[4] NETTRAN_DUMMY_4985 NETTRAN_DUMMY_4986 
+ NETTRAN_DUMMY_4987 DFF_X1 
Xdata_out_reg_5_ n1126 n82_G2B1I2 data_out[5] NETTRAN_DUMMY_4988 NETTRAN_DUMMY_4989 
+ NETTRAN_DUMMY_4990 DFF_X1 
Xdata_out_reg_6_ n1118 n82_G2B1I2 n2026 NETTRAN_DUMMY_4991 NETTRAN_DUMMY_4992 NETTRAN_DUMMY_4993 DFF_X1 
Xdata_out_reg_7_ n1117 n82_G2B1I7 data_out[7] NETTRAN_DUMMY_4994 NETTRAN_DUMMY_4995 
+ NETTRAN_DUMMY_4996 DFF_X1 
Xdata_out_reg_8_ n554 n125_G2B1I5 data_out[8] NETTRAN_DUMMY_4997 NETTRAN_DUMMY_4998 
+ NETTRAN_DUMMY_4999 DFF_X1 
Xdata_out_reg_9_ n553 n125_G2B1I5 data_out[9] NETTRAN_DUMMY_5000 NETTRAN_DUMMY_5001 
+ NETTRAN_DUMMY_5002 DFF_X1 
Xdata_out_reg_10_ n1098 n82_G2B1I8 data_out[10] NETTRAN_DUMMY_5003 NETTRAN_DUMMY_5004 
+ NETTRAN_DUMMY_5005 DFF_X1 
Xdata_out_reg_11_ n1093 n82_G2B1I2 data_out[11] NETTRAN_DUMMY_5006 NETTRAN_DUMMY_5007 
+ NETTRAN_DUMMY_5008 DFF_X1 
Xdata_out_reg_12_ n1092 n125 data_out[12] NETTRAN_DUMMY_5009 NETTRAN_DUMMY_5010 
+ NETTRAN_DUMMY_5011 DFF_X1 
Xdata_out_reg_13_ n1086 n125 data_out[13] NETTRAN_DUMMY_5012 NETTRAN_DUMMY_5013 
+ NETTRAN_DUMMY_5014 DFF_X1 
Xdata_out_reg_14_ n1082 n125 n2024 NETTRAN_DUMMY_5015 NETTRAN_DUMMY_5016 NETTRAN_DUMMY_5017 DFF_X1 
Xdata_out_reg_15_ n1076 n125 data_out[15] NETTRAN_DUMMY_5018 NETTRAN_DUMMY_5019 
+ NETTRAN_DUMMY_5020 DFF_X1 
Xdata_out_reg_16_ n2028 n125_G2B1I5 data_out[16] NETTRAN_DUMMY_5021 NETTRAN_DUMMY_5022 
+ NETTRAN_DUMMY_5023 DFF_X1 
Xdata_out_reg_17_ n1066 n125_G2B1I5 data_out[17] NETTRAN_DUMMY_5024 NETTRAN_DUMMY_5025 
+ NETTRAN_DUMMY_5026 DFF_X1 
Xdata_out_reg_18_ n1065 n125_G2B1I1 data_out[18] NETTRAN_DUMMY_5027 NETTRAN_DUMMY_5028 
+ NETTRAN_DUMMY_5029 DFF_X1 
Xdata_out_reg_19_ n1056 n125_G2B1I1 data_out[19] NETTRAN_DUMMY_5030 NETTRAN_DUMMY_5031 
+ NETTRAN_DUMMY_5032 DFF_X1 
Xdata_out_reg_20_ n1051 n125_G2B1I1 data_out[20] NETTRAN_DUMMY_5033 NETTRAN_DUMMY_5034 
+ NETTRAN_DUMMY_5035 DFF_X1 
Xdata_out_reg_21_ n2030 n125_G2B1I3 data_out[21] NETTRAN_DUMMY_5036 NETTRAN_DUMMY_5037 
+ NETTRAN_DUMMY_5038 DFF_X1 
Xdata_out_reg_22_ n1044 n125_G2B1I6 data_out[22] NETTRAN_DUMMY_5039 NETTRAN_DUMMY_5040 
+ NETTRAN_DUMMY_5041 DFF_X1 
Xdata_out_reg_23_ n1035 n125_G2B1I1 data_out[23] NETTRAN_DUMMY_5042 NETTRAN_DUMMY_5043 
+ NETTRAN_DUMMY_5044 DFF_X1 
Xdata_out_reg_24_ n1029 n125_G2B1I6 data_out[24] NETTRAN_DUMMY_5045 NETTRAN_DUMMY_5046 
+ NETTRAN_DUMMY_5047 DFF_X1 
Xdata_out_reg_25_ n1023 n76 data_out[25] NETTRAN_DUMMY_5048 NETTRAN_DUMMY_5049 NETTRAN_DUMMY_5050 DFF_X1 
Xdata_out_reg_26_ n552 n125_G2B1I3 data_out[26] NETTRAN_DUMMY_5051 NETTRAN_DUMMY_5052 
+ NETTRAN_DUMMY_5053 DFF_X1 
Xdata_out_reg_27_ n309 n125_G2B1I1 data_out[27] NETTRAN_DUMMY_5054 NETTRAN_DUMMY_5055 
+ NETTRAN_DUMMY_5056 DFF_X1 
Xdata_out_reg_28_ n1009 n76 data_out[28] NETTRAN_DUMMY_5057 NETTRAN_DUMMY_5058 NETTRAN_DUMMY_5059 DFF_X1 
Xdata_out_reg_29_ n1003 n125_G2B1I6 data_out[29] NETTRAN_DUMMY_5060 NETTRAN_DUMMY_5061 
+ NETTRAN_DUMMY_5062 DFF_X1 
Xdata_out_reg_30_ n997 n125_G2B1I6 data_out[30] NETTRAN_DUMMY_5063 NETTRAN_DUMMY_5064 
+ NETTRAN_DUMMY_5065 DFF_X1 
Xdata_out_reg_31_ n308 n125_G2B1I6 data_out[31] NETTRAN_DUMMY_5066 NETTRAN_DUMMY_5067 
+ NETTRAN_DUMMY_5068 DFF_X1 
Xdata_out_reg_32_ n985 n78_G2B1I4 data_out[32] NETTRAN_DUMMY_5069 NETTRAN_DUMMY_5070 
+ NETTRAN_DUMMY_5071 DFF_X1 
Xdata_out_reg_33_ n979 n78_G2B1I4 data_out[33] NETTRAN_DUMMY_5072 NETTRAN_DUMMY_5073 
+ NETTRAN_DUMMY_5074 DFF_X1 
Xdata_out_reg_34_ n973 n78 data_out[34] NETTRAN_DUMMY_5075 NETTRAN_DUMMY_5076 NETTRAN_DUMMY_5077 DFF_X1 
Xdata_out_reg_35_ n968 n78_G2B1I6 data_out[35] NETTRAN_DUMMY_5078 NETTRAN_DUMMY_5079 
+ NETTRAN_DUMMY_5080 DFF_X1 
Xdata_out_reg_36_ n962 n78_G2B1I1 data_out[36] NETTRAN_DUMMY_5081 NETTRAN_DUMMY_5082 
+ NETTRAN_DUMMY_5083 DFF_X1 
Xdata_out_reg_37_ n956 n78_G2B1I1 data_out[37] NETTRAN_DUMMY_5084 NETTRAN_DUMMY_5085 
+ NETTRAN_DUMMY_5086 DFF_X1 
Xdata_out_reg_38_ n950 n78_G2B1I5 data_out[38] NETTRAN_DUMMY_5087 NETTRAN_DUMMY_5088 
+ NETTRAN_DUMMY_5089 DFF_X1 
Xdata_out_reg_39_ n944 n78_G2B1I4 data_out[39] NETTRAN_DUMMY_5090 NETTRAN_DUMMY_5091 
+ NETTRAN_DUMMY_5092 DFF_X1 
Xdata_out_reg_40_ n942 n78 data_out[40] NETTRAN_DUMMY_5093 NETTRAN_DUMMY_5094 NETTRAN_DUMMY_5095 DFF_X1 
Xdata_out_reg_41_ n936 n78 data_out[41] NETTRAN_DUMMY_5096 NETTRAN_DUMMY_5097 NETTRAN_DUMMY_5098 DFF_X1 
Xdata_out_reg_42_ n573 n78_G2B1I5 data_out[42] NETTRAN_DUMMY_5099 NETTRAN_DUMMY_5100 
+ NETTRAN_DUMMY_5101 DFF_X1 
Xdata_out_reg_43_ n924 n78_G2B1I5 data_out[43] NETTRAN_DUMMY_5102 NETTRAN_DUMMY_5103 
+ NETTRAN_DUMMY_5104 DFF_X1 
Xdata_out_reg_44_ n918 n78_G2B1I1 data_out[44] NETTRAN_DUMMY_5105 NETTRAN_DUMMY_5106 
+ NETTRAN_DUMMY_5107 DFF_X1 
Xdata_out_reg_45_ n307 n78_G2B1I1 data_out[45] NETTRAN_DUMMY_5108 NETTRAN_DUMMY_5109 
+ NETTRAN_DUMMY_5110 DFF_X1 
Xdata_out_reg_46_ n906 n78_G2B1I5 data_out[46] NETTRAN_DUMMY_5111 NETTRAN_DUMMY_5112 
+ NETTRAN_DUMMY_5113 DFF_X1 
Xdata_out_reg_47_ n900 n78_G2B1I1 data_out[47] NETTRAN_DUMMY_5114 NETTRAN_DUMMY_5115 
+ NETTRAN_DUMMY_5116 DFF_X1 
Xdata_out_reg_48_ n894 n125_G2B1I1 data_out[48] NETTRAN_DUMMY_5117 NETTRAN_DUMMY_5118 
+ NETTRAN_DUMMY_5119 DFF_X1 
Xdata_out_reg_49_ n888 n125_G2B1I4 data_out[49] NETTRAN_DUMMY_5120 NETTRAN_DUMMY_5121 
+ NETTRAN_DUMMY_5122 DFF_X1 
Xdata_out_reg_50_ n882 n125_G2B1I3 data_out[50] NETTRAN_DUMMY_5123 NETTRAN_DUMMY_5124 
+ NETTRAN_DUMMY_5125 DFF_X1 
Xdata_out_reg_51_ n306 n125_G2B1I3 data_out[51] NETTRAN_DUMMY_5126 NETTRAN_DUMMY_5127 
+ NETTRAN_DUMMY_5128 DFF_X1 
Xdata_out_reg_52_ n870 n125_G2B1I6 data_out[52] NETTRAN_DUMMY_5129 NETTRAN_DUMMY_5130 
+ NETTRAN_DUMMY_5131 DFF_X1 
Xdata_out_reg_53_ n864 n125_G2B1I6 data_out[53] NETTRAN_DUMMY_5132 NETTRAN_DUMMY_5133 
+ NETTRAN_DUMMY_5134 DFF_X1 
Xdata_out_reg_54_ n858 n125_G2B1I6 data_out[54] NETTRAN_DUMMY_5135 NETTRAN_DUMMY_5136 
+ NETTRAN_DUMMY_5137 DFF_X1 
Xdata_out_reg_55_ n852 n125_G2B1I1 data_out[55] NETTRAN_DUMMY_5138 NETTRAN_DUMMY_5139 
+ NETTRAN_DUMMY_5140 DFF_X1 
Xdata_out_reg_56_ n846 n125_G2B1I4 data_out[56] NETTRAN_DUMMY_5141 NETTRAN_DUMMY_5142 
+ NETTRAN_DUMMY_5143 DFF_X1 
Xdata_out_reg_57_ n305 n125_G2B1I4 data_out[57] NETTRAN_DUMMY_5144 NETTRAN_DUMMY_5145 
+ NETTRAN_DUMMY_5146 DFF_X1 
Xdata_out_reg_58_ n836 n125_G2B1I5 data_out[58] NETTRAN_DUMMY_5147 NETTRAN_DUMMY_5148 
+ NETTRAN_DUMMY_5149 DFF_X1 
Xdata_out_reg_59_ n2029 n125_G2B1I5 data_out[59] NETTRAN_DUMMY_5150 NETTRAN_DUMMY_5151 
+ NETTRAN_DUMMY_5152 DFF_X1 
Xdata_out_reg_60_ n824 n125_G2B1I5 data_out[60] NETTRAN_DUMMY_5153 NETTRAN_DUMMY_5154 
+ NETTRAN_DUMMY_5155 DFF_X1 
Xdata_out_reg_61_ n818 n125_G2B1I5 data_out[61] NETTRAN_DUMMY_5156 NETTRAN_DUMMY_5157 
+ NETTRAN_DUMMY_5158 DFF_X1 
Xdata_out_reg_62_ n2027 n125_G2B1I4 data_out[62] NETTRAN_DUMMY_5159 NETTRAN_DUMMY_5160 
+ NETTRAN_DUMMY_5161 DFF_X1 
Xdata_out_reg_63_ n304 n125_G2B1I4 data_out[63] NETTRAN_DUMMY_5162 NETTRAN_DUMMY_5163 
+ NETTRAN_DUMMY_5164 DFF_X1 
Xvalid_out_reg n256 n76_G2B1I3 valid_out NETTRAN_DUMMY_5165 NETTRAN_DUMMY_5166 NETTRAN_DUMMY_5167 DFF_X1 
Xz2_reg_51_ n571 n80_G2B1I4 NETTRAN_DUMMY_5168 n139 NETTRAN_DUMMY_5169 NETTRAN_DUMMY_5170 DFF_X1 
Xz2_reg_38_ n570 n80_G2B1I6 z2_next[51] n152 NETTRAN_DUMMY_5171 NETTRAN_DUMMY_5172 DFF_X1 
Xz2_reg_25_ n567 n80 z2_next[38] n165 NETTRAN_DUMMY_5173 NETTRAN_DUMMY_5174 DFF_X1 
Xz2_reg_12_ n565 n80 z2_next[25] n178 NETTRAN_DUMMY_5175 NETTRAN_DUMMY_5176 DFF_X1 
Xz2_reg_57_ n564 n80_G2B1I6 NETTRAN_DUMMY_5177 n133 NETTRAN_DUMMY_5178 NETTRAN_DUMMY_5179 DFF_X1 
Xz2_reg_44_ n563 n84_G2B1I2 z2_next[57] n146 NETTRAN_DUMMY_5180 NETTRAN_DUMMY_5181 DFF_X1 
Xz2_reg_31_ n561 n84_G2B1I2 z2_next[44] n159 NETTRAN_DUMMY_5182 NETTRAN_DUMMY_5183 DFF_X1 
Xz2_reg_18_ n765 n76_G2B1I4 z2_next[31] n172 NETTRAN_DUMMY_5184 NETTRAN_DUMMY_5185 DFF_X1 
Xz2_reg_63_ n560 n76_G2B1I4 z2[63] n124 NETTRAN_DUMMY_5186 NETTRAN_DUMMY_5187 DFF_X1 
Xz2_reg_50_ n559 n76_G2B1I1 z2_next[63] n140 NETTRAN_DUMMY_5188 NETTRAN_DUMMY_5189 DFF_X1 
Xz2_reg_37_ n558 n84_G2B1I2 z2_next[50] n153 NETTRAN_DUMMY_5190 NETTRAN_DUMMY_5191 DFF_X1 
XU76 IN0 n254 n50 n261 n43 n539 NETTRAN_DUMMY_5192 NETTRAN_DUMMY_5193 OAI221_X1 
XU75 IN0 n255 n53 n260 n46 n542 NETTRAN_DUMMY_5194 NETTRAN_DUMMY_5195 OAI221_X1 
XU74 IN0 n254 n729 n261 n24 n520 NETTRAN_DUMMY_5196 NETTRAN_DUMMY_5197 OAI221_X1 
XU73 IN2 n255 n1646 n258 n41 n537 NETTRAN_DUMMY_5198 NETTRAN_DUMMY_5199 OAI221_X1 
XU72 IN0 n254 n20 n261 n13 n509 NETTRAN_DUMMY_5200 NETTRAN_DUMMY_5201 OAI221_X1 
XU71 rstn n254 n13 n261 n1676 n502 NETTRAN_DUMMY_5202 NETTRAN_DUMMY_5203 OAI221_X1 
XU70 rstn n254 n16 n261 n9 n505 NETTRAN_DUMMY_5204 NETTRAN_DUMMY_5205 OAI221_X1 
XU69 IN0 n254 n9 n261 n1719 n498 NETTRAN_DUMMY_5206 NETTRAN_DUMMY_5207 OAI221_X1 
XU68 IN2 n255 n698 n258 n1729 n543 NETTRAN_DUMMY_5208 NETTRAN_DUMMY_5209 OAI221_X1 
XU67 IN0 n254 n703 n261 n12 n508 NETTRAN_DUMMY_5210 NETTRAN_DUMMY_5211 OAI221_X1 
XU66 IN0 n254 n12 n261 n5 n501 NETTRAN_DUMMY_5212 NETTRAN_DUMMY_5213 OAI221_X1 
XU65 rstn n254 n29 n258 n22 n518 NETTRAN_DUMMY_5214 NETTRAN_DUMMY_5215 OAI221_X1 
XU64 IN2 n255 n22 n258 n1797 n511 NETTRAN_DUMMY_5216 NETTRAN_DUMMY_5217 OAI221_X1 
XU63 IN0 n254 n1797 n258 n806 n504 NETTRAN_DUMMY_5218 NETTRAN_DUMMY_5219 OAI221_X1 
XU62 IN2 n255 n806 n260 n1 n497 NETTRAN_DUMMY_5220 NETTRAN_DUMMY_5221 OAI221_X1 
XU61 IN0 n254 n11 n261 n4 n500 NETTRAN_DUMMY_5222 NETTRAN_DUMMY_5223 OAI221_X1 
XU60 IN2 n255 n719 n258 n42 n538 NETTRAN_DUMMY_5224 NETTRAN_DUMMY_5225 OAI221_X1 
XU59 IN0 n254 n14 n261 n1881 n503 NETTRAN_DUMMY_5226 NETTRAN_DUMMY_5227 OAI221_X1 
XU58 IN0 n254 n1886 n261 n726 n541 NETTRAN_DUMMY_5228 NETTRAN_DUMMY_5229 OAI221_X1 
XU57 rstn n254 n732 n261 n10 n506 NETTRAN_DUMMY_5230 NETTRAN_DUMMY_5231 OAI221_X1 
XU56 IN0 n254 n10 n261 n3 n499 NETTRAN_DUMMY_5232 NETTRAN_DUMMY_5233 OAI221_X1 
XU55 IN3 n2531 n735 n260 n1931 n472 NETTRAN_DUMMY_5234 NETTRAN_DUMMY_5235 OAI221_X1 
XU54 IN3 n2531 n109 n260 n85 n458 NETTRAN_DUMMY_5236 NETTRAN_DUMMY_5237 OAI221_X1 
XU53 IN2 n255 n119 n260 n95 n468 NETTRAN_DUMMY_5238 NETTRAN_DUMMY_5239 OAI221_X1 
XU52 IN2 n255 n120 n260 n96 n469 NETTRAN_DUMMY_5240 NETTRAN_DUMMY_5241 OAI221_X1 
XU51 IN3 n2531 n96 n259 n67 n445 NETTRAN_DUMMY_5242 NETTRAN_DUMMY_5243 OAI221_X1 
XU50 IN3 n2531 n121 n260 n97 n470 NETTRAN_DUMMY_5244 NETTRAN_DUMMY_5245 OAI221_X1 
XU49 IN3 n2531 n122 n259 n98 n471 NETTRAN_DUMMY_5246 NETTRAN_DUMMY_5247 OAI221_X1 
XU48 IN3 n2531 n118 n260 n94 n467 NETTRAN_DUMMY_5248 NETTRAN_DUMMY_5249 OAI221_X1 
XU47 IN3 n2531 n94 n260 n65 n443 NETTRAN_DUMMY_5250 NETTRAN_DUMMY_5251 OAI221_X1 
XU46 IN3 n2531 n597 n259 n90 n463 NETTRAN_DUMMY_5252 NETTRAN_DUMMY_5253 OAI221_X1 
XU45 IN3 n2531 n115 n259 n91 n464 NETTRAN_DUMMY_5254 NETTRAN_DUMMY_5255 OAI221_X1 
XU44 IN3 n2531 n110 n260 n86 n459 NETTRAN_DUMMY_5256 NETTRAN_DUMMY_5257 OAI221_X1 
XU43 IN3 n2531 n609 n259 n1300 n465 NETTRAN_DUMMY_5258 NETTRAN_DUMMY_5259 OAI221_X1 
XU42 IN3 n2531 n111 n259 n87 n460 NETTRAN_DUMMY_5260 NETTRAN_DUMMY_5261 OAI221_X1 
XU41 IN3 n2531 n117 n259 n93 n466 NETTRAN_DUMMY_5262 NETTRAN_DUMMY_5263 OAI221_X1 
XU40 IN3 n2531 n112 n259 n88 n461 NETTRAN_DUMMY_5264 NETTRAN_DUMMY_5265 OAI221_X1 
XU39 IN3 n2531 n113 n259 n89 n462 NETTRAN_DUMMY_5266 NETTRAN_DUMMY_5267 OAI221_X1 
XU38 IN2 n255 n140 n258 n124 n376 NETTRAN_DUMMY_5268 NETTRAN_DUMMY_5269 OAI221_X1 
XU37 n252 n1080 N2610 NETTRAN_DUMMY_5270 NETTRAN_DUMMY_5271 NOR2_X1 
XU36 n252 n331 N2600 NETTRAN_DUMMY_5272 NETTRAN_DUMMY_5273 NOR2_X1 
XU35 n252 n333 N2590 NETTRAN_DUMMY_5274 NETTRAN_DUMMY_5275 NOR2_X1 
XU34 n252 n1090 N2580 NETTRAN_DUMMY_5276 NETTRAN_DUMMY_5277 NOR2_X1 
XU33 n252 n1095 N2570 NETTRAN_DUMMY_5278 NETTRAN_DUMMY_5279 NOR2_X1 
XU32 n252 n1100 N2560 NETTRAN_DUMMY_5280 NETTRAN_DUMMY_5281 NOR2_X1 
XU31 n252 n1105 N2550 NETTRAN_DUMMY_5282 NETTRAN_DUMMY_5283 NOR2_X1 
XU19 IN0 n255 n188 NETTRAN_DUMMY_5284 NETTRAN_DUMMY_5285 NAND2_X1 
XU18 n188 n258 NETTRAN_DUMMY_5286 NETTRAN_DUMMY_5287 BUF_X2 
XU17 n187 n257 NETTRAN_DUMMY_5288 NETTRAN_DUMMY_5289 BUF_X2 
XU15 n187 n255 NETTRAN_DUMMY_5290 NETTRAN_DUMMY_5291 BUF_X2 
XU14 n187 n254 NETTRAN_DUMMY_5292 NETTRAN_DUMMY_5293 BUF_X2 
XU13 n187 n2531 NETTRAN_DUMMY_5294 NETTRAN_DUMMY_5295 BUF_X2 
XU441 n373 n374 n372 NETTRAN_DUMMY_5296 NETTRAN_DUMMY_5297 XOR2_X1 
XU440 n369 n370 n368 NETTRAN_DUMMY_5298 NETTRAN_DUMMY_5299 XOR2_X1 
XU439 n365 n366 n364 NETTRAN_DUMMY_5300 NETTRAN_DUMMY_5301 XOR2_X1 
XU438 n361 n362 n360 NETTRAN_DUMMY_5302 NETTRAN_DUMMY_5303 XOR2_X1 
XU437 n357 n358 n356 NETTRAN_DUMMY_5304 NETTRAN_DUMMY_5305 XOR2_X1 
XU436 n353 n354 n352 NETTRAN_DUMMY_5306 NETTRAN_DUMMY_5307 XOR2_X1 
XU435 n83 z1[45] n220 NETTRAN_DUMMY_5308 NETTRAN_DUMMY_5309 XOR2_X1 
XU434 n201 n220 n351 NETTRAN_DUMMY_5310 NETTRAN_DUMMY_5311 XOR2_X1 
XU433 n350 n351 n349 NETTRAN_DUMMY_5312 NETTRAN_DUMMY_5313 XOR2_X1 
XU432 n81 z1[46] n219 NETTRAN_DUMMY_5314 NETTRAN_DUMMY_5315 XOR2_X1 
XU431 n200 n219 n348 NETTRAN_DUMMY_5316 NETTRAN_DUMMY_5317 XOR2_X1 
XU430 n347 n348 n346 NETTRAN_DUMMY_5318 NETTRAN_DUMMY_5319 XOR2_X1 
XU429 n79 z1[47] n218 NETTRAN_DUMMY_5320 NETTRAN_DUMMY_5321 XOR2_X1 
XU428 n199 n218 n345 NETTRAN_DUMMY_5322 NETTRAN_DUMMY_5323 XOR2_X1 
XU427 n344 n345 n343 NETTRAN_DUMMY_5324 NETTRAN_DUMMY_5325 XOR2_X1 
XU426 n77 z1[48] n217 NETTRAN_DUMMY_5326 NETTRAN_DUMMY_5327 XOR2_X1 
XU425 n198 n217 n342 NETTRAN_DUMMY_5328 NETTRAN_DUMMY_5329 XOR2_X1 
XU424 n232 n342 n341 NETTRAN_DUMMY_5330 NETTRAN_DUMMY_5331 XOR2_X1 
XU423 n75 z1[49] n216 NETTRAN_DUMMY_5332 NETTRAN_DUMMY_5333 XOR2_X1 
XU169 IN2 n255 n161 n258 n1573 n397 NETTRAN_DUMMY_5334 NETTRAN_DUMMY_5335 OAI221_X1 
XU168 IN2 n255 n1573 n258 n135 n384 NETTRAN_DUMMY_5336 NETTRAN_DUMMY_5337 OAI221_X1 
XU167 IN2 n255 n167 n258 n154 n403 NETTRAN_DUMMY_5338 NETTRAN_DUMMY_5339 OAI221_X1 
XU166 IN2 n255 n141 n258 n126 n377 NETTRAN_DUMMY_5340 NETTRAN_DUMMY_5341 OAI221_X1 
XU165 IN2 n255 n173 n258 n160 n409 NETTRAN_DUMMY_5342 NETTRAN_DUMMY_5343 OAI221_X1 
XU164 IN2 n255 n160 n258 n147 n396 NETTRAN_DUMMY_5344 NETTRAN_DUMMY_5345 OAI221_X1 
XU163 IN2 n255 n147 n258 n134 n383 NETTRAN_DUMMY_5346 NETTRAN_DUMMY_5347 OAI221_X1 
XU162 IN0 n255 n166 n260 n153 n402 NETTRAN_DUMMY_5348 NETTRAN_DUMMY_5349 OAI221_X1 
XU161 IN2 n255 n153 n140 n258 n389 NETTRAN_DUMMY_5350 NETTRAN_DUMMY_5351 OAI221_X1 
XU160 IN0 n255 n172 n260 n774 n408 NETTRAN_DUMMY_5352 NETTRAN_DUMMY_5353 OAI221_X1 
XU159 IN0 n255 n774 n260 n146 n395 NETTRAN_DUMMY_5354 NETTRAN_DUMMY_5355 OAI221_X1 
XU158 IN0 n257 n146 n261 n133 n382 NETTRAN_DUMMY_5356 NETTRAN_DUMMY_5357 OAI221_X1 
XU157 IN0 n257 n165 n261 n152 n401 NETTRAN_DUMMY_5358 NETTRAN_DUMMY_5359 OAI221_X1 
XU156 IN0 n257 n152 n261 n139 n388 NETTRAN_DUMMY_5360 NETTRAN_DUMMY_5361 OAI221_X1 
XU155 n225 n623 NETTRAN_DUMMY_5362 NETTRAN_DUMMY_5363 INV_X1 
XU154 IN3 n623 n2531 n259 n735 n496 NETTRAN_DUMMY_5364 NETTRAN_DUMMY_5365 OAI221_X1 
XU153 IN2 n231 n255 n258 n698 n550 NETTRAN_DUMMY_5366 NETTRAN_DUMMY_5367 OAI221_X1 
XU152 IN2 n226 n255 n258 n719 n545 NETTRAN_DUMMY_5368 NETTRAN_DUMMY_5369 OAI221_X1 
XU151 IN0 n229 n254 n261 n1886 n548 NETTRAN_DUMMY_5370 NETTRAN_DUMMY_5371 OAI221_X1 
XU150 n221 n619 NETTRAN_DUMMY_5372 NETTRAN_DUMMY_5373 INV_X1 
XU149 IN2 n619 n255 n260 n119 n492 NETTRAN_DUMMY_5374 NETTRAN_DUMMY_5375 OAI221_X1 
XU148 n224 n622 NETTRAN_DUMMY_5376 NETTRAN_DUMMY_5377 INV_X1 
XU147 IN3 n622 n2531 n259 n122 n495 NETTRAN_DUMMY_5378 NETTRAN_DUMMY_5379 OAI221_X1 
XU146 IN3 n206 n2531 n259 n104 n477 NETTRAN_DUMMY_5380 NETTRAN_DUMMY_5381 OAI221_X1 
XU145 IN2 n202 n255 n260 n100 n473 NETTRAN_DUMMY_5382 NETTRAN_DUMMY_5383 OAI221_X1 
XU144 IN3 n203 n2531 n259 n101 n474 NETTRAN_DUMMY_5384 NETTRAN_DUMMY_5385 OAI221_X1 
XU143 IN3 n218 n2531 n259 n609 n489 NETTRAN_DUMMY_5386 NETTRAN_DUMMY_5387 OAI221_X1 
XU142 IN3 n204 n2531 n259 n102 n475 NETTRAN_DUMMY_5388 NETTRAN_DUMMY_5389 OAI221_X1 
XU141 IN0 n200 n257 n259 n183 n432 NETTRAN_DUMMY_5390 NETTRAN_DUMMY_5391 OAI221_X1 
XU140 rstn n198 n254 n258 n667 n430 NETTRAN_DUMMY_5392 NETTRAN_DUMMY_5393 OAI221_X1 
XU139 IN2 n197 n255 n258 n1581 n429 NETTRAN_DUMMY_5394 NETTRAN_DUMMY_5395 OAI221_X1 
XU138 n261 n27 n254 n34 n523 NETTRAN_DUMMY_5396 NETTRAN_DUMMY_5397 OAI22_X1 
XU137 n261 n30 n254 n37 n526 NETTRAN_DUMMY_5398 NETTRAN_DUMMY_5399 OAI22_X1 
XU136 n261 n23 n254 n30 n519 NETTRAN_DUMMY_5400 NETTRAN_DUMMY_5401 OAI22_X1 
XU135 n261 n700 n254 n40 n529 NETTRAN_DUMMY_5402 NETTRAN_DUMMY_5403 OAI22_X1 
XU134 n261 n701 n254 n700 n522 NETTRAN_DUMMY_5404 NETTRAN_DUMMY_5405 OAI22_X1 
XU133 n261 n29 n254 n36 n525 NETTRAN_DUMMY_5406 NETTRAN_DUMMY_5407 OAI22_X1 
XU132 n260 n32 n257 n39 n528 NETTRAN_DUMMY_5408 NETTRAN_DUMMY_5409 OAI22_X1 
XU131 n260 n25 n2531 n32 n521 NETTRAN_DUMMY_5410 NETTRAN_DUMMY_5411 OAI22_X1 
XU130 n260 n18 n2531 n25 n514 NETTRAN_DUMMY_5412 NETTRAN_DUMMY_5413 OAI22_X1 
XU129 n260 n28 n255 n35 n524 NETTRAN_DUMMY_5414 NETTRAN_DUMMY_5415 OAI22_X1 
XU128 n258 n21 n254 n28 n517 NETTRAN_DUMMY_5416 NETTRAN_DUMMY_5417 OAI22_X1 
XU127 n261 n729 n254 n727 n527 NETTRAN_DUMMY_5418 NETTRAN_DUMMY_5419 OAI22_X1 
XU126 n260 n70 n2531 n99 n448 NETTRAN_DUMMY_5420 NETTRAN_DUMMY_5421 OAI22_X1 
XU125 n260 n56 n2531 n85 n434 NETTRAN_DUMMY_5422 NETTRAN_DUMMY_5423 OAI22_X1 
XU124 n260 n66 n255 n95 n444 NETTRAN_DUMMY_5424 NETTRAN_DUMMY_5425 OAI22_X1 
XU123 n260 n77 n255 n105 n454 NETTRAN_DUMMY_5426 NETTRAN_DUMMY_5427 OAI22_X1 
XU122 n259 n79 n2531 n2001 n455 NETTRAN_DUMMY_5428 NETTRAN_DUMMY_5429 OAI22_X1 
XU121 n259 n68 n2531 n97 n446 NETTRAN_DUMMY_5430 NETTRAN_DUMMY_5431 OAI22_X1 
XU120 n259 n81 n257 n107 n456 NETTRAN_DUMMY_5432 NETTRAN_DUMMY_5433 OAI22_X1 
XU119 n259 n69 n257 n98 n447 NETTRAN_DUMMY_5434 NETTRAN_DUMMY_5435 OAI22_X1 
XU118 n259 n83 n257 n108 n457 NETTRAN_DUMMY_5436 NETTRAN_DUMMY_5437 OAI22_X1 
XU117 n260 n75 n2531 n104 n453 NETTRAN_DUMMY_5438 NETTRAN_DUMMY_5439 OAI22_X1 
XU116 n260 n71 n255 n100 n449 NETTRAN_DUMMY_5440 NETTRAN_DUMMY_5441 OAI22_X1 
XU115 n259 n62 n2531 n91 n440 NETTRAN_DUMMY_5442 NETTRAN_DUMMY_5443 OAI22_X1 
XU114 n259 n72 n2531 n101 n450 NETTRAN_DUMMY_5444 NETTRAN_DUMMY_5445 OAI22_X1 
XU113 n259 n58 n2531 n87 n436 NETTRAN_DUMMY_5446 NETTRAN_DUMMY_5447 OAI22_X1 
XU112 n259 n73 n2531 n102 n451 NETTRAN_DUMMY_5448 NETTRAN_DUMMY_5449 OAI22_X1 
XU111 n259 n59 n257 n88 n437 NETTRAN_DUMMY_5450 NETTRAN_DUMMY_5451 OAI22_X1 
XU110 n259 n74 n257 n103 n452 NETTRAN_DUMMY_5452 NETTRAN_DUMMY_5453 OAI22_X1 
XU109 n259 n60 n2531 n89 n438 NETTRAN_DUMMY_5454 NETTRAN_DUMMY_5455 OAI22_X1 
XU108 n259 n1396 n257 n184 n420 NETTRAN_DUMMY_5456 NETTRAN_DUMMY_5457 OAI22_X1 
XU107 n260 n1152 n257 n1418 n413 NETTRAN_DUMMY_5458 NETTRAN_DUMMY_5459 OAI22_X1 
XU106 n259 n170 n257 n183 n419 NETTRAN_DUMMY_5460 NETTRAN_DUMMY_5461 OAI22_X1 
XU105 n259 n1491 n257 n182 n418 NETTRAN_DUMMY_5462 NETTRAN_DUMMY_5463 OAI22_X1 
XU104 n258 n1537 n254 n667 n417 NETTRAN_DUMMY_5464 NETTRAN_DUMMY_5465 OAI22_X1 
XU103 n258 n161 n255 n174 n410 NETTRAN_DUMMY_5466 NETTRAN_DUMMY_5467 OAI22_X1 
XU102 n258 n167 n255 n1581 n416 NETTRAN_DUMMY_5468 NETTRAN_DUMMY_5469 OAI22_X1 
XU101 n258 n166 n254 n179 n415 NETTRAN_DUMMY_5470 NETTRAN_DUMMY_5471 OAI22_X1 
XU100 n259 n165 n257 n178 n414 NETTRAN_DUMMY_5472 NETTRAN_DUMMY_5473 OAI22_X1 
XU99 n258 n1646 n255 n1640 n544 NETTRAN_DUMMY_5474 NETTRAN_DUMMY_5475 OAI22_X1 
XU98 n258 n34 n254 n41 n530 NETTRAN_DUMMY_5476 NETTRAN_DUMMY_5477 OAI22_X1 
XU97 n261 n37 n254 n44 n533 NETTRAN_DUMMY_5478 NETTRAN_DUMMY_5479 OAI22_X1 
XU96 n258 n40 n255 n47 n536 NETTRAN_DUMMY_5480 NETTRAN_DUMMY_5481 OAI22_X1 
XU95 n261 n36 n254 n43 n532 NETTRAN_DUMMY_5482 NETTRAN_DUMMY_5483 OAI22_X1 
XU94 n260 n39 n257 n46 n535 NETTRAN_DUMMY_5484 NETTRAN_DUMMY_5485 OAI22_X1 
XU93 n260 n11 n257 n18 n507 NETTRAN_DUMMY_5486 NETTRAN_DUMMY_5487 OAI22_X1 
XU92 n258 n35 n255 n42 n531 NETTRAN_DUMMY_5488 NETTRAN_DUMMY_5489 OAI22_X1 
XU91 n261 n727 n257 n726 n534 NETTRAN_DUMMY_5490 NETTRAN_DUMMY_5491 OAI22_X1 
XU90 n261 n144 n257 n157 n393 NETTRAN_DUMMY_5492 NETTRAN_DUMMY_5493 OAI22_X1 
XU89 n258 n142 n254 n155 n391 NETTRAN_DUMMY_5494 NETTRAN_DUMMY_5495 OAI22_X1 
XU88 n258 n141 n255 n154 n390 NETTRAN_DUMMY_5496 NETTRAN_DUMMY_5497 OAI22_X1 
XU87 n222 n620 NETTRAN_DUMMY_5498 NETTRAN_DUMMY_5499 INV_X1 
XU86 IN2 n620 n255 n260 n120 n493 NETTRAN_DUMMY_5500 NETTRAN_DUMMY_5501 OAI221_X1 
XU85 n223 n621 NETTRAN_DUMMY_5502 NETTRAN_DUMMY_5503 INV_X1 
XU84 IN3 n621 n2531 n260 n121 n494 NETTRAN_DUMMY_5504 NETTRAN_DUMMY_5505 OAI221_X1 
XU83 IN3 n220 n2531 n260 n118 n491 NETTRAN_DUMMY_5506 NETTRAN_DUMMY_5507 OAI221_X1 
XU82 IN3 n216 n2531 n259 n597 n487 NETTRAN_DUMMY_5508 NETTRAN_DUMMY_5509 OAI221_X1 
XU81 IN3 n219 n2531 n259 n117 n490 NETTRAN_DUMMY_5510 NETTRAN_DUMMY_5511 OAI221_X1 
XU80 IN3 n205 n257 n259 n103 n476 NETTRAN_DUMMY_5512 NETTRAN_DUMMY_5513 OAI221_X1 
XU79 IN0 n254 n27 n261 n20 n516 NETTRAN_DUMMY_5514 NETTRAN_DUMMY_5515 OAI221_X1 
XU78 IN0 n254 n51 n261 n44 n540 NETTRAN_DUMMY_5516 NETTRAN_DUMMY_5517 OAI221_X1 
XU77 IN0 n254 n701 n261 n703 n515 NETTRAN_DUMMY_5518 NETTRAN_DUMMY_5519 OAI221_X1 
XU262 z2_next[20] z3_next[20] n320 NETTRAN_DUMMY_5520 NETTRAN_DUMMY_5521 XNOR2_X1 
XU261 n320 n206 n319 NETTRAN_DUMMY_5522 NETTRAN_DUMMY_5523 XNOR2_X1 
XU260 n185 n1053 N266 NETTRAN_DUMMY_5524 NETTRAN_DUMMY_5525 NOR2_X1 
XU259 z2_next[19] z3_next[19] n322 NETTRAN_DUMMY_5526 NETTRAN_DUMMY_5527 XNOR2_X1 
XU258 n322 n207 n321 NETTRAN_DUMMY_5528 NETTRAN_DUMMY_5529 XNOR2_X1 
XU257 n185 n1058 N265 NETTRAN_DUMMY_5530 NETTRAN_DUMMY_5531 NOR2_X1 
XU256 z3_next[18] n189 n324 NETTRAN_DUMMY_5532 NETTRAN_DUMMY_5533 XNOR2_X1 
XU255 n324 n208 n323 NETTRAN_DUMMY_5534 NETTRAN_DUMMY_5535 XNOR2_X1 
XU254 n185 n1063 N264 NETTRAN_DUMMY_5536 NETTRAN_DUMMY_5537 NOR2_X1 
XU253 z3_next[17] n190 n326 NETTRAN_DUMMY_5538 NETTRAN_DUMMY_5539 XNOR2_X1 
XU252 n326 n209 n325 NETTRAN_DUMMY_5540 NETTRAN_DUMMY_5541 XNOR2_X1 
XU251 n252 n1068 N263 NETTRAN_DUMMY_5542 NETTRAN_DUMMY_5543 NOR2_X1 
XU250 z3_next[16] n191 n328 NETTRAN_DUMMY_5544 NETTRAN_DUMMY_5545 XNOR2_X1 
XU249 n328 n210 n327 NETTRAN_DUMMY_5546 NETTRAN_DUMMY_5547 XNOR2_X1 
XU248 n252 n1073 N262 NETTRAN_DUMMY_5548 NETTRAN_DUMMY_5549 NOR2_X1 
XU247 z3_next[39] z3_next[63] n344 NETTRAN_DUMMY_5550 NETTRAN_DUMMY_5551 XNOR2_X1 
XU246 n252 n1110 N2540 NETTRAN_DUMMY_5552 NETTRAN_DUMMY_5553 NOR2_X1 
XU245 z3_next[38] z3_next[62] n347 NETTRAN_DUMMY_5554 NETTRAN_DUMMY_5555 XNOR2_X1 
XU244 n252 n1115 N253 NETTRAN_DUMMY_5556 NETTRAN_DUMMY_5557 NOR2_X1 
XU243 z3_next[37] z3_next[61] n350 NETTRAN_DUMMY_5558 NETTRAN_DUMMY_5559 XNOR2_X1 
XU242 n252 n1120 N2520 NETTRAN_DUMMY_5560 NETTRAN_DUMMY_5561 NOR2_X1 
XU241 n140 n355 n354 NETTRAN_DUMMY_5562 NETTRAN_DUMMY_5563 XNOR2_X1 
XU240 z2_next[44] n221 n353 NETTRAN_DUMMY_5564 NETTRAN_DUMMY_5565 XNOR2_X1 
XU239 n252 n1124 N251 NETTRAN_DUMMY_5566 NETTRAN_DUMMY_5567 NOR2_X1 
XU238 n141 n359 n358 NETTRAN_DUMMY_5568 NETTRAN_DUMMY_5569 XNOR2_X1 
XU237 z2_next[43] n222 n357 NETTRAN_DUMMY_5570 NETTRAN_DUMMY_5571 XNOR2_X1 
XU236 n252 n1129 N2500 NETTRAN_DUMMY_5572 NETTRAN_DUMMY_5573 NOR2_X1 
XU235 z2_next[42] n223 n361 NETTRAN_DUMMY_5574 NETTRAN_DUMMY_5575 XNOR2_X1 
XU234 n142 n363 n362 NETTRAN_DUMMY_5576 NETTRAN_DUMMY_5577 XNOR2_X1 
XU233 n252 n1134 N249 NETTRAN_DUMMY_5578 NETTRAN_DUMMY_5579 NOR2_X1 
XU232 n143 n367 n366 NETTRAN_DUMMY_5580 NETTRAN_DUMMY_5581 XNOR2_X1 
XU231 z2_next[41] n224 n365 NETTRAN_DUMMY_5582 NETTRAN_DUMMY_5583 XNOR2_X1 
XU230 n250 n1139 N2480 NETTRAN_DUMMY_5584 NETTRAN_DUMMY_5585 NOR2_X1 
XU229 n144 n371 n370 NETTRAN_DUMMY_5586 NETTRAN_DUMMY_5587 XNOR2_X1 
XU228 z2_next[40] n225 n369 NETTRAN_DUMMY_5588 NETTRAN_DUMMY_5589 XNOR2_X1 
XU227 n246 n1144 N247 NETTRAN_DUMMY_5590 NETTRAN_DUMMY_5591 NOR2_X1 
XU226 n1152 n375 n374 NETTRAN_DUMMY_5592 NETTRAN_DUMMY_5593 XNOR2_X1 
XU225 n576 n244 n373 NETTRAN_DUMMY_5594 NETTRAN_DUMMY_5595 XNOR2_X1 
XU224 n185 n1148 N2460 NETTRAN_DUMMY_5596 NETTRAN_DUMMY_5597 NOR2_X1 
XU222 n261 n732 n254 n24 n513 NETTRAN_DUMMY_5598 NETTRAN_DUMMY_5599 OAI22_X1 
XU221 n261 n16 n254 n23 n512 NETTRAN_DUMMY_5600 NETTRAN_DUMMY_5601 OAI22_X1 
XU220 n261 n14 n254 n21 n510 NETTRAN_DUMMY_5602 NETTRAN_DUMMY_5603 OAI22_X1 
XU219 ce IN3 n187 NETTRAN_DUMMY_5604 NETTRAN_DUMMY_5605 NAND2_X1 
XU218 n258 n1640 n232 n255 n551 NETTRAN_DUMMY_5606 NETTRAN_DUMMY_5607 OAI22_X1 
XU217 n261 n1681 n228 n254 n547 NETTRAN_DUMMY_5608 NETTRAN_DUMMY_5609 OAI22_X1 
XU216 n261 n1765 n227 n254 n546 NETTRAN_DUMMY_5610 NETTRAN_DUMMY_5611 OAI22_X1 
XU215 n260 n53 n230 n255 n549 NETTRAN_DUMMY_5612 NETTRAN_DUMMY_5613 OAI22_X1 
XU214 n259 n2001 n208 n2531 n479 NETTRAN_DUMMY_5614 NETTRAN_DUMMY_5615 OAI22_X1 
XU213 n259 n107 n209 n2531 n480 NETTRAN_DUMMY_5616 NETTRAN_DUMMY_5617 OAI22_X1 
XU212 n259 n587 n210 n257 n481 NETTRAN_DUMMY_5618 NETTRAN_DUMMY_5619 OAI22_X1 
XU211 n259 n115 n217 n2531 n488 NETTRAN_DUMMY_5620 NETTRAN_DUMMY_5621 OAI22_X1 
XU210 n260 n110 n212 n2531 n483 NETTRAN_DUMMY_5622 NETTRAN_DUMMY_5623 OAI22_X1 
XU209 n261 n1418 n194 n257 n426 NETTRAN_DUMMY_5624 NETTRAN_DUMMY_5625 OAI22_X1 
XU208 n261 n176 n193 n257 n425 NETTRAN_DUMMY_5626 NETTRAN_DUMMY_5627 OAI22_X1 
XU207 n191 n624 NETTRAN_DUMMY_5628 NETTRAN_DUMMY_5629 INV_X1 
XU206 n258 n174 n624 n255 n423 NETTRAN_DUMMY_5630 NETTRAN_DUMMY_5631 OAI22_X1 
XU205 n260 n109 n211 n2531 n482 NETTRAN_DUMMY_5632 NETTRAN_DUMMY_5633 OAI22_X1 
XU204 n260 n105 n207 n255 n478 NETTRAN_DUMMY_5634 NETTRAN_DUMMY_5635 OAI22_X1 
XU203 n259 n111 n213 n2531 n484 NETTRAN_DUMMY_5636 NETTRAN_DUMMY_5637 OAI22_X1 
XU202 n259 n112 n214 n2531 n485 NETTRAN_DUMMY_5638 NETTRAN_DUMMY_5639 OAI22_X1 
XU201 n259 n113 n215 n257 n486 NETTRAN_DUMMY_5640 NETTRAN_DUMMY_5641 OAI22_X1 
XU200 n259 n184 n201 n257 n433 NETTRAN_DUMMY_5642 NETTRAN_DUMMY_5643 OAI22_X1 
XU199 n259 n182 n199 n257 n431 NETTRAN_DUMMY_5644 NETTRAN_DUMMY_5645 OAI22_X1 
XU198 n258 n175 n192 n254 n424 NETTRAN_DUMMY_5646 NETTRAN_DUMMY_5647 OAI22_X1 
XU197 n190 n625 NETTRAN_DUMMY_5648 NETTRAN_DUMMY_5649 INV_X1 
XU196 n258 n173 n625 n255 n422 NETTRAN_DUMMY_5650 NETTRAN_DUMMY_5651 OAI22_X1 
XU195 n258 n179 n196 n254 n428 NETTRAN_DUMMY_5652 NETTRAN_DUMMY_5653 OAI22_X1 
XU194 n189 n626 NETTRAN_DUMMY_5654 NETTRAN_DUMMY_5655 INV_X1 
XU193 n260 n172 n626 n255 n421 NETTRAN_DUMMY_5656 NETTRAN_DUMMY_5657 OAI22_X1 
XU192 n261 n178 n195 n257 n427 NETTRAN_DUMMY_5658 NETTRAN_DUMMY_5659 OAI22_X1 
XU191 IN3 n2531 n90 n260 n1974 n439 NETTRAN_DUMMY_5660 NETTRAN_DUMMY_5661 OAI221_X1 
XU190 IN3 n2531 n86 n260 n57 n435 NETTRAN_DUMMY_5662 NETTRAN_DUMMY_5663 OAI221_X1 
XU189 IN3 n2531 n1300 n259 n63 n441 NETTRAN_DUMMY_5664 NETTRAN_DUMMY_5665 OAI221_X1 
XU188 IN3 n2531 n93 n259 n64 n442 NETTRAN_DUMMY_5666 NETTRAN_DUMMY_5667 OAI221_X1 
XU187 IN3 n257 n1396 n259 n643 n407 NETTRAN_DUMMY_5668 NETTRAN_DUMMY_5669 OAI221_X1 
XU186 IN0 n257 n643 n259 n1406 n394 NETTRAN_DUMMY_5670 NETTRAN_DUMMY_5671 OAI221_X1 
XU185 IN0 n257 n1406 n261 n132 n381 NETTRAN_DUMMY_5672 NETTRAN_DUMMY_5673 OAI221_X1 
XU184 IN0 n257 n1152 n261 n151 n400 NETTRAN_DUMMY_5674 NETTRAN_DUMMY_5675 OAI221_X1 
XU183 IN0 n257 n151 n261 n138 n387 NETTRAN_DUMMY_5676 NETTRAN_DUMMY_5677 OAI221_X1 
XU182 IN3 n257 n170 n259 n157 n406 NETTRAN_DUMMY_5678 NETTRAN_DUMMY_5679 OAI221_X1 
XU181 IN0 n257 n144 n261 n131 n380 NETTRAN_DUMMY_5680 NETTRAN_DUMMY_5681 OAI221_X1 
XU180 IN0 n257 n176 n259 n1470 n412 NETTRAN_DUMMY_5682 NETTRAN_DUMMY_5683 OAI221_X1 
XU179 IN0 n257 n1470 n259 n150 n399 NETTRAN_DUMMY_5684 NETTRAN_DUMMY_5685 OAI221_X1 
XU178 IN0 n257 n150 n261 n137 n386 NETTRAN_DUMMY_5686 NETTRAN_DUMMY_5687 OAI221_X1 
XU177 IN3 n257 n1491 n259 n156 n405 NETTRAN_DUMMY_5688 NETTRAN_DUMMY_5689 OAI221_X1 
XU176 IN0 n257 n156 n261 n143 n392 NETTRAN_DUMMY_5690 NETTRAN_DUMMY_5691 OAI221_X1 
XU175 IN0 n254 n143 n261 n130 n379 NETTRAN_DUMMY_5692 NETTRAN_DUMMY_5693 OAI221_X1 
XU174 rstn n254 n175 n258 n162 n411 NETTRAN_DUMMY_5694 NETTRAN_DUMMY_5695 OAI221_X1 
XU173 rstn n254 n162 n258 n149 n398 NETTRAN_DUMMY_5696 NETTRAN_DUMMY_5697 OAI221_X1 
XU172 rstn n254 n149 n258 n136 n385 NETTRAN_DUMMY_5698 NETTRAN_DUMMY_5699 OAI221_X1 
XU171 rstn n254 n1537 n258 n155 n404 NETTRAN_DUMMY_5700 NETTRAN_DUMMY_5701 OAI221_X1 
XU170 rstn n254 n142 n258 n128 n378 NETTRAN_DUMMY_5702 NETTRAN_DUMMY_5703 OAI221_X1 
XU355 n20 z2_next[51] n25800 NETTRAN_DUMMY_5704 NETTRAN_DUMMY_5705 XNOR2_X1 
XU354 z1_next[51] n25800 n25700 NETTRAN_DUMMY_5706 NETTRAN_DUMMY_5707 XNOR2_X1 
XU353 n185 n878 N297 NETTRAN_DUMMY_5708 NETTRAN_DUMMY_5709 NOR2_X1 
XU352 n21 z2_next[50] n26000 NETTRAN_DUMMY_5710 NETTRAN_DUMMY_5711 XNOR2_X1 
XU351 z1_next[50] n26000 n25900 NETTRAN_DUMMY_5712 NETTRAN_DUMMY_5713 XNOR2_X1 
XU350 n252 n886 N296 NETTRAN_DUMMY_5714 NETTRAN_DUMMY_5715 NOR2_X1 
XU349 n22 z2_next[49] n2620 NETTRAN_DUMMY_5716 NETTRAN_DUMMY_5717 XNOR2_X1 
XU348 z1_next[49] n2620 n26100 NETTRAN_DUMMY_5718 NETTRAN_DUMMY_5719 XNOR2_X1 
XU347 n185 n890 N295 NETTRAN_DUMMY_5720 NETTRAN_DUMMY_5721 NOR2_X1 
XU346 n23 z2_next[48] n2640 NETTRAN_DUMMY_5722 NETTRAN_DUMMY_5723 XNOR2_X1 
XU345 z1_next[48] n2640 n2630 NETTRAN_DUMMY_5724 NETTRAN_DUMMY_5725 XNOR2_X1 
XU344 n185 n896 N294 NETTRAN_DUMMY_5726 NETTRAN_DUMMY_5727 NOR2_X1 
XU343 n24 z2_next[47] n2660 NETTRAN_DUMMY_5728 NETTRAN_DUMMY_5729 XNOR2_X1 
XU342 z1_next[47] n2660 n2650 NETTRAN_DUMMY_5730 NETTRAN_DUMMY_5731 XNOR2_X1 
XU341 n248 n902 N293 NETTRAN_DUMMY_5732 NETTRAN_DUMMY_5733 NOR2_X1 
XU340 n25 z2_next[46] n2680 NETTRAN_DUMMY_5734 NETTRAN_DUMMY_5735 XNOR2_X1 
XU339 z1_next[46] n2680 n2670 NETTRAN_DUMMY_5736 NETTRAN_DUMMY_5737 XNOR2_X1 
XU338 n248 n908 N292 NETTRAN_DUMMY_5738 NETTRAN_DUMMY_5739 NOR2_X1 
XU337 n26 z2_next[45] n2700 NETTRAN_DUMMY_5740 NETTRAN_DUMMY_5741 XNOR2_X1 
XU336 z1_next[45] n2700 n2690 NETTRAN_DUMMY_5742 NETTRAN_DUMMY_5743 XNOR2_X1 
XU335 n246 n914 N291 NETTRAN_DUMMY_5744 NETTRAN_DUMMY_5745 NOR2_X1 
XU334 n27 z2_next[44] n2720 NETTRAN_DUMMY_5746 NETTRAN_DUMMY_5747 XNOR2_X1 
XU333 z1_next[44] n2720 n2710 NETTRAN_DUMMY_5748 NETTRAN_DUMMY_5749 XNOR2_X1 
XU332 n246 n920 N290 NETTRAN_DUMMY_5750 NETTRAN_DUMMY_5751 NOR2_X1 
XU331 n28 z2_next[43] n2740 NETTRAN_DUMMY_5752 NETTRAN_DUMMY_5753 XNOR2_X1 
XU330 z1_next[43] n2740 n2730 NETTRAN_DUMMY_5754 NETTRAN_DUMMY_5755 XNOR2_X1 
XU329 n246 n926 N289 NETTRAN_DUMMY_5756 NETTRAN_DUMMY_5757 NOR2_X1 
XU328 n29 z2_next[42] n2760 NETTRAN_DUMMY_5758 NETTRAN_DUMMY_5759 XNOR2_X1 
XU327 z1_next[42] n2760 n2750 NETTRAN_DUMMY_5760 NETTRAN_DUMMY_5761 XNOR2_X1 
XU326 n246 n932 N288 NETTRAN_DUMMY_5762 NETTRAN_DUMMY_5763 NOR2_X1 
XU325 n30 z2_next[41] n2780 NETTRAN_DUMMY_5764 NETTRAN_DUMMY_5765 XNOR2_X1 
XU324 z1_next[41] n2780 n2770 NETTRAN_DUMMY_5766 NETTRAN_DUMMY_5767 XNOR2_X1 
XU323 n246 n938 N287 NETTRAN_DUMMY_5768 NETTRAN_DUMMY_5769 NOR2_X1 
XU322 n31 z2_next[40] n2800 NETTRAN_DUMMY_5770 NETTRAN_DUMMY_5771 XNOR2_X1 
XU321 z1_next[40] n2800 n2790 NETTRAN_DUMMY_5772 NETTRAN_DUMMY_5773 XNOR2_X1 
XU320 n246 n940 N286 NETTRAN_DUMMY_5774 NETTRAN_DUMMY_5775 NOR2_X1 
XU319 n32 z2_next[39] n2820 NETTRAN_DUMMY_5776 NETTRAN_DUMMY_5777 XNOR2_X1 
XU318 z1_next[39] n2820 n2810 NETTRAN_DUMMY_5778 NETTRAN_DUMMY_5779 XNOR2_X1 
XU317 n246 n946 N285 NETTRAN_DUMMY_5780 NETTRAN_DUMMY_5781 NOR2_X1 
XU316 n33 z2_next[38] n2840 NETTRAN_DUMMY_5782 NETTRAN_DUMMY_5783 XNOR2_X1 
XU315 z1_next[38] n2840 n2830 NETTRAN_DUMMY_5784 NETTRAN_DUMMY_5785 XNOR2_X1 
XU314 n246 n952 N284 NETTRAN_DUMMY_5786 NETTRAN_DUMMY_5787 NOR2_X1 
XU313 n34 z2_next[37] n2860 NETTRAN_DUMMY_5788 NETTRAN_DUMMY_5789 XNOR2_X1 
XU312 z1_next[37] n2860 n2850 NETTRAN_DUMMY_5790 NETTRAN_DUMMY_5791 XNOR2_X1 
XU311 n246 n958 N283 NETTRAN_DUMMY_5792 NETTRAN_DUMMY_5793 NOR2_X1 
XU310 n35 z2_next[36] n2880 NETTRAN_DUMMY_5794 NETTRAN_DUMMY_5795 XNOR2_X1 
XU309 z1_next[36] n2880 n2870 NETTRAN_DUMMY_5796 NETTRAN_DUMMY_5797 XNOR2_X1 
XU308 n246 n964 N282 NETTRAN_DUMMY_5798 NETTRAN_DUMMY_5799 NOR2_X1 
XU307 n36 z2_next[35] n2900 NETTRAN_DUMMY_5800 NETTRAN_DUMMY_5801 XNOR2_X1 
XU306 z1_next[35] n2900 n2890 NETTRAN_DUMMY_5802 NETTRAN_DUMMY_5803 XNOR2_X1 
XU305 n246 n970 N281 NETTRAN_DUMMY_5804 NETTRAN_DUMMY_5805 NOR2_X1 
XU304 n37 z2_next[34] n2920 NETTRAN_DUMMY_5806 NETTRAN_DUMMY_5807 XNOR2_X1 
XU303 z1_next[34] n2920 n2910 NETTRAN_DUMMY_5808 NETTRAN_DUMMY_5809 XNOR2_X1 
XU302 n246 n977 N280 NETTRAN_DUMMY_5810 NETTRAN_DUMMY_5811 NOR2_X1 
XU301 n38 z2_next[33] n2940 NETTRAN_DUMMY_5812 NETTRAN_DUMMY_5813 XNOR2_X1 
XU300 z1_next[33] n2940 n2930 NETTRAN_DUMMY_5814 NETTRAN_DUMMY_5815 XNOR2_X1 
XU299 n246 n981 N279 NETTRAN_DUMMY_5816 NETTRAN_DUMMY_5817 NOR2_X1 
XU298 n39 z2_next[32] n2960 NETTRAN_DUMMY_5818 NETTRAN_DUMMY_5819 XNOR2_X1 
XU297 z1_next[32] n2960 n2950 NETTRAN_DUMMY_5820 NETTRAN_DUMMY_5821 XNOR2_X1 
XU296 n246 n987 N278 NETTRAN_DUMMY_5822 NETTRAN_DUMMY_5823 NOR2_X1 
XU295 n40 z2_next[31] n2980 NETTRAN_DUMMY_5824 NETTRAN_DUMMY_5825 XNOR2_X1 
XU294 z1_next[31] n2980 n2970 NETTRAN_DUMMY_5826 NETTRAN_DUMMY_5827 XNOR2_X1 
XU293 n185 n993 N277 NETTRAN_DUMMY_5828 NETTRAN_DUMMY_5829 NOR2_X1 
XU292 n41 z2_next[30] n3000 NETTRAN_DUMMY_5830 NETTRAN_DUMMY_5831 XNOR2_X1 
XU291 z1_next[30] n3000 n2990 NETTRAN_DUMMY_5832 NETTRAN_DUMMY_5833 XNOR2_X1 
XU290 n185 n999 N276 NETTRAN_DUMMY_5834 NETTRAN_DUMMY_5835 NOR2_X1 
XU289 n42 z2_next[29] n3020 NETTRAN_DUMMY_5836 NETTRAN_DUMMY_5837 XNOR2_X1 
XU288 z1_next[29] n3020 n3010 NETTRAN_DUMMY_5838 NETTRAN_DUMMY_5839 XNOR2_X1 
XU287 n185 n1007 N275 NETTRAN_DUMMY_5840 NETTRAN_DUMMY_5841 NOR2_X1 
XU286 n43 z2_next[28] n3040 NETTRAN_DUMMY_5842 NETTRAN_DUMMY_5843 XNOR2_X1 
XU285 z1_next[28] n3040 n3030 NETTRAN_DUMMY_5844 NETTRAN_DUMMY_5845 XNOR2_X1 
XU284 n185 n1011 N274 NETTRAN_DUMMY_5846 NETTRAN_DUMMY_5847 NOR2_X1 
XU283 n44 z2_next[27] n3060 NETTRAN_DUMMY_5848 NETTRAN_DUMMY_5849 XNOR2_X1 
XU282 z1_next[27] n3060 n3050 NETTRAN_DUMMY_5850 NETTRAN_DUMMY_5851 XNOR2_X1 
XU281 n185 n1016 N273 NETTRAN_DUMMY_5852 NETTRAN_DUMMY_5853 NOR2_X1 
XU280 n45 z2_next[26] n3080 NETTRAN_DUMMY_5854 NETTRAN_DUMMY_5855 XNOR2_X1 
XU279 z1_next[26] n3080 n3070 NETTRAN_DUMMY_5856 NETTRAN_DUMMY_5857 XNOR2_X1 
XU278 n185 n1020 N272 NETTRAN_DUMMY_5858 NETTRAN_DUMMY_5859 NOR2_X1 
XU277 n46 z2_next[25] n310 NETTRAN_DUMMY_5860 NETTRAN_DUMMY_5861 XNOR2_X1 
XU276 z1_next[25] n310 n3090 NETTRAN_DUMMY_5862 NETTRAN_DUMMY_5863 XNOR2_X1 
XU275 n185 n1025 N271 NETTRAN_DUMMY_5864 NETTRAN_DUMMY_5865 NOR2_X1 
XU274 z2_next[24] z3_next[24] n312 NETTRAN_DUMMY_5866 NETTRAN_DUMMY_5867 XNOR2_X1 
XU273 n312 n202 n311 NETTRAN_DUMMY_5868 NETTRAN_DUMMY_5869 XNOR2_X1 
XU272 n185 n1031 N270 NETTRAN_DUMMY_5870 NETTRAN_DUMMY_5871 NOR2_X1 
XU271 z2_next[23] z3_next[23] n314 NETTRAN_DUMMY_5872 NETTRAN_DUMMY_5873 XNOR2_X1 
XU270 n314 n203 n313 NETTRAN_DUMMY_5874 NETTRAN_DUMMY_5875 XNOR2_X1 
XU269 n185 n1037 N269 NETTRAN_DUMMY_5876 NETTRAN_DUMMY_5877 NOR2_X1 
XU268 z2_next[22] z3_next[22] n316 NETTRAN_DUMMY_5878 NETTRAN_DUMMY_5879 XNOR2_X1 
XU267 n316 n204 n315 NETTRAN_DUMMY_5880 NETTRAN_DUMMY_5881 XNOR2_X1 
XU266 n185 n1042 N268 NETTRAN_DUMMY_5882 NETTRAN_DUMMY_5883 NOR2_X1 
XU265 z2_next[21] z3_next[21] n318 NETTRAN_DUMMY_5884 NETTRAN_DUMMY_5885 XNOR2_X1 
XU264 n318 n205 n317 NETTRAN_DUMMY_5886 NETTRAN_DUMMY_5887 XNOR2_X1 
XU263 n185 n1047 N267 NETTRAN_DUMMY_5888 NETTRAN_DUMMY_5889 NOR2_X1 
XU467 n13 z3_next[34] n363 NETTRAN_DUMMY_5890 NETTRAN_DUMMY_5891 XNOR2_X1 
XU466 n12 z3_next[35] n359 NETTRAN_DUMMY_5892 NETTRAN_DUMMY_5893 XNOR2_X1 
XU465 n1797 z3_next[32] n371 NETTRAN_DUMMY_5894 NETTRAN_DUMMY_5895 XNOR2_X1 
XU464 n11 z3_next[36] n355 NETTRAN_DUMMY_5896 NETTRAN_DUMMY_5897 XNOR2_X1 
XU463 n14 z3_next[33] n367 NETTRAN_DUMMY_5898 NETTRAN_DUMMY_5899 XNOR2_X1 
XU462 n16 z3_next[31] n375 NETTRAN_DUMMY_5900 NETTRAN_DUMMY_5901 XNOR2_X1 
XU461 z3[62] z3_next[45] n227 NETTRAN_DUMMY_5902 NETTRAN_DUMMY_5903 XNOR2_X1 
XU460 z3[61] z3_next[44] n228 NETTRAN_DUMMY_5904 NETTRAN_DUMMY_5905 XNOR2_X1 
XU459 z3[59] z3_next[42] n230 NETTRAN_DUMMY_5906 NETTRAN_DUMMY_5907 XNOR2_X1 
XU458 z3[57] z3_next[40] n232 NETTRAN_DUMMY_5908 NETTRAN_DUMMY_5909 XNOR2_X1 
XU457 n130 n149 n192 NETTRAN_DUMMY_5910 NETTRAN_DUMMY_5911 XNOR2_X1 
XU456 n131 n150 n193 NETTRAN_DUMMY_5912 NETTRAN_DUMMY_5913 XNOR2_X1 
XU455 n132 n151 n194 NETTRAN_DUMMY_5914 NETTRAN_DUMMY_5915 XNOR2_X1 
XU454 n133 n152 n195 NETTRAN_DUMMY_5916 NETTRAN_DUMMY_5917 XNOR2_X1 
XU453 n134 n153 n196 NETTRAN_DUMMY_5918 NETTRAN_DUMMY_5919 XNOR2_X1 
XU452 n137 n156 n199 NETTRAN_DUMMY_5920 NETTRAN_DUMMY_5921 XNOR2_X1 
XU451 n139 n158 n201 NETTRAN_DUMMY_5922 NETTRAN_DUMMY_5923 XNOR2_X1 
XU450 z3[63] z3_next[46] n226 NETTRAN_DUMMY_5924 NETTRAN_DUMMY_5925 XNOR2_X1 
XU449 z3[60] z3_next[43] n229 NETTRAN_DUMMY_5926 NETTRAN_DUMMY_5927 XNOR2_X1 
XU448 z3[58] z3_next[41] n231 NETTRAN_DUMMY_5928 NETTRAN_DUMMY_5929 XNOR2_X1 
XU447 n135 n154 n197 NETTRAN_DUMMY_5930 NETTRAN_DUMMY_5931 XNOR2_X1 
XU446 n136 n155 n198 NETTRAN_DUMMY_5932 NETTRAN_DUMMY_5933 XNOR2_X1 
XU445 n138 n157 n200 NETTRAN_DUMMY_5934 NETTRAN_DUMMY_5935 XNOR2_X1 
XU444 n66 n1974 n207 NETTRAN_DUMMY_5936 NETTRAN_DUMMY_5937 XNOR2_X1 
XU443 n68 n63 n209 NETTRAN_DUMMY_5938 NETTRAN_DUMMY_5939 XNOR2_X1 
XU442 n69 n64 n210 NETTRAN_DUMMY_5940 NETTRAN_DUMMY_5941 XNOR2_X1 
XU405 n67 n62 n208 NETTRAN_DUMMY_5942 NETTRAN_DUMMY_5943 XNOR2_X1 
XU404 z2[63] n146 n189 NETTRAN_DUMMY_5944 NETTRAN_DUMMY_5945 XNOR2_X1 
XU403 z2[62] n147 n190 NETTRAN_DUMMY_5946 NETTRAN_DUMMY_5947 XNOR2_X1 
XU402 z2[61] n1573 n191 NETTRAN_DUMMY_5948 NETTRAN_DUMMY_5949 XNOR2_X1 
XU401 z1[43] n86 n222 NETTRAN_DUMMY_5950 NETTRAN_DUMMY_5951 XNOR2_X1 
XU400 z1[44] n85 n221 NETTRAN_DUMMY_5952 NETTRAN_DUMMY_5953 XNOR2_X1 
XU399 z1[42] n87 n223 NETTRAN_DUMMY_5954 NETTRAN_DUMMY_5955 XNOR2_X1 
XU398 z1[41] n88 n224 NETTRAN_DUMMY_5956 NETTRAN_DUMMY_5957 XNOR2_X1 
XU397 z1[40] n89 n225 NETTRAN_DUMMY_5958 NETTRAN_DUMMY_5959 XNOR2_X1 
XU396 n65 n60 n206 NETTRAN_DUMMY_5960 NETTRAN_DUMMY_5961 XNOR2_X1 
XU395 n1974 n56 n202 NETTRAN_DUMMY_5962 NETTRAN_DUMMY_5963 XNOR2_X1 
XU394 n63 n58 n204 NETTRAN_DUMMY_5964 NETTRAN_DUMMY_5965 XNOR2_X1 
XU393 n64 n59 n205 NETTRAN_DUMMY_5966 NETTRAN_DUMMY_5967 XNOR2_X1 
XU392 n62 n57 n203 NETTRAN_DUMMY_5968 NETTRAN_DUMMY_5969 XNOR2_X1 
XU391 n90 z2_next[58] n244 NETTRAN_DUMMY_5970 NETTRAN_DUMMY_5971 XNOR2_X1 
XU390 n806 z2_next[63] n234 NETTRAN_DUMMY_5972 NETTRAN_DUMMY_5973 XNOR2_X1 
XU389 n576 n234 n233 NETTRAN_DUMMY_5974 NETTRAN_DUMMY_5975 XNOR2_X1 
XU388 n252 n808 N3091 NETTRAN_DUMMY_5976 NETTRAN_DUMMY_5977 NOR2_X1 
XU387 n9 z2_next[62] n236 NETTRAN_DUMMY_5978 NETTRAN_DUMMY_5979 XNOR2_X1 
XU386 z1_next[62] n236 n235 NETTRAN_DUMMY_5980 NETTRAN_DUMMY_5981 XNOR2_X1 
XU385 n252 n814 N3081 NETTRAN_DUMMY_5982 NETTRAN_DUMMY_5983 NOR2_X1 
XU384 n10 z2_next[61] n238 NETTRAN_DUMMY_5984 NETTRAN_DUMMY_5985 XNOR2_X1 
XU383 z1_next[61] n238 n237 NETTRAN_DUMMY_5986 NETTRAN_DUMMY_5987 XNOR2_X1 
XU382 n252 n820 N3071 NETTRAN_DUMMY_5988 NETTRAN_DUMMY_5989 NOR2_X1 
XU381 n11 z2_next[60] n240 NETTRAN_DUMMY_5990 NETTRAN_DUMMY_5991 XNOR2_X1 
XU380 z1_next[60] n240 n239 NETTRAN_DUMMY_5992 NETTRAN_DUMMY_5993 XNOR2_X1 
XU379 n252 n826 N3061 NETTRAN_DUMMY_5994 NETTRAN_DUMMY_5995 NOR2_X1 
XU378 n12 z2_next[59] n242 NETTRAN_DUMMY_5996 NETTRAN_DUMMY_5997 XNOR2_X1 
XU377 z1_next[59] n242 n241 NETTRAN_DUMMY_5998 NETTRAN_DUMMY_5999 XNOR2_X1 
XU376 n252 n832 N3051 NETTRAN_DUMMY_6000 NETTRAN_DUMMY_6001 NOR2_X1 
XU375 z3_next[58] n244 n243 NETTRAN_DUMMY_6002 NETTRAN_DUMMY_6003 XNOR2_X1 
XU374 n252 n838 N3041 NETTRAN_DUMMY_6004 NETTRAN_DUMMY_6005 NOR2_X1 
XU373 n14 z2_next[57] n24600 NETTRAN_DUMMY_6006 NETTRAN_DUMMY_6007 XNOR2_X1 
XU372 z1_next[57] n24600 n245 NETTRAN_DUMMY_6008 NETTRAN_DUMMY_6009 XNOR2_X1 
XU371 n185 n843 N303 NETTRAN_DUMMY_6010 NETTRAN_DUMMY_6011 NOR2_X1 
XU370 n1797 z2_next[56] n24800 NETTRAN_DUMMY_6012 NETTRAN_DUMMY_6013 XNOR2_X1 
XU369 z1_next[56] n24800 n2470 NETTRAN_DUMMY_6014 NETTRAN_DUMMY_6015 XNOR2_X1 
XU368 n185 n848 N302 NETTRAN_DUMMY_6016 NETTRAN_DUMMY_6017 NOR2_X1 
XU367 n16 z2_next[55] n25000 NETTRAN_DUMMY_6018 NETTRAN_DUMMY_6019 XNOR2_X1 
XU366 z1_next[55] n25000 n2490 NETTRAN_DUMMY_6020 NETTRAN_DUMMY_6021 XNOR2_X1 
XU365 n185 n854 N301 NETTRAN_DUMMY_6022 NETTRAN_DUMMY_6023 NOR2_X1 
XU364 n17 z2_next[54] n25200 NETTRAN_DUMMY_6024 NETTRAN_DUMMY_6025 XNOR2_X1 
XU363 z1_next[54] n25200 n2510 NETTRAN_DUMMY_6026 NETTRAN_DUMMY_6027 XNOR2_X1 
XU362 n185 n860 N300 NETTRAN_DUMMY_6028 NETTRAN_DUMMY_6029 NOR2_X1 
XU361 n18 z2_next[53] n25400 NETTRAN_DUMMY_6030 NETTRAN_DUMMY_6031 XNOR2_X1 
XU360 z1_next[53] n25400 n2530 NETTRAN_DUMMY_6032 NETTRAN_DUMMY_6033 XNOR2_X1 
XU359 n185 n868 N299 NETTRAN_DUMMY_6034 NETTRAN_DUMMY_6035 NOR2_X1 
XU358 n19 z2_next[52] n25600 NETTRAN_DUMMY_6036 NETTRAN_DUMMY_6037 XNOR2_X1 
XU357 z1_next[52] n25600 n25500 NETTRAN_DUMMY_6038 NETTRAN_DUMMY_6039 XNOR2_X1 
XU356 n185 n874 N298 NETTRAN_DUMMY_6040 NETTRAN_DUMMY_6041 NOR2_X1 
XCLKBUF_X1_G2B1I1 n78 n78_G2B1I1 NETTRAN_DUMMY_6042 NETTRAN_DUMMY_6043 CLKBUF_X1 
XCLKBUF_X1_G2B1I2 n78 n78_G2B1I2 NETTRAN_DUMMY_6044 NETTRAN_DUMMY_6045 CLKBUF_X1 
XCLKBUF_X1_G2B1I4 n78 n78_G2B1I4 NETTRAN_DUMMY_6046 NETTRAN_DUMMY_6047 CLKBUF_X1 
XCLKBUF_X1_G2B1I5 n78 n78_G2B1I5 NETTRAN_DUMMY_6048 NETTRAN_DUMMY_6049 CLKBUF_X1 
XCLKBUF_X1_G2B1I6 n78 n78_G2B1I6 NETTRAN_DUMMY_6050 NETTRAN_DUMMY_6051 CLKBUF_X1 
XCLKBUF_X1_G2B1I7 n78 n78_G2B1I7 NETTRAN_DUMMY_6052 NETTRAN_DUMMY_6053 CLKBUF_X1 
XCLKBUF_X1_G2B1I8 n78 n78_G2B1I8 NETTRAN_DUMMY_6054 NETTRAN_DUMMY_6055 CLKBUF_X1 
XCLKBUF_X1_G2B1I11 n125 n125_G2B1I1 NETTRAN_DUMMY_6056 NETTRAN_DUMMY_6057 CLKBUF_X1 
XCLKBUF_X1_G2B1I31 n125 n125_G2B1I3 NETTRAN_DUMMY_6058 NETTRAN_DUMMY_6059 CLKBUF_X1 
XCLKBUF_X1_G2B1I41 n125 n125_G2B1I4 NETTRAN_DUMMY_6060 NETTRAN_DUMMY_6061 CLKBUF_X1 
XCLKBUF_X1_G2B1I51 n125 n125_G2B1I5 NETTRAN_DUMMY_6062 NETTRAN_DUMMY_6063 CLKBUF_X1 
XCLKBUF_X1_G2B1I61 n125 n125_G2B1I6 NETTRAN_DUMMY_6064 NETTRAN_DUMMY_6065 CLKBUF_X1 
XCLKBUF_X1_G2B1I22 n84 n84_G2B1I2 NETTRAN_DUMMY_6066 NETTRAN_DUMMY_6067 CLKBUF_X1 
XCLKBUF_X1_G2B1I32 n84 n84_G2B1I3 NETTRAN_DUMMY_6068 NETTRAN_DUMMY_6069 CLKBUF_X1 
XCLKBUF_X1_G2B1I42 n84 n84_G2B1I4 NETTRAN_DUMMY_6070 NETTRAN_DUMMY_6071 CLKBUF_X1 
XCLKBUF_X1_G2B1I52 n84 n84_G2B1I5 NETTRAN_DUMMY_6072 NETTRAN_DUMMY_6073 CLKBUF_X1 
XCLKBUF_X1_G2B1I62 n84 n84_G2B1I6 NETTRAN_DUMMY_6074 NETTRAN_DUMMY_6075 CLKBUF_X1 
XCLKBUF_X1_G2B1I13 n76 n76_G2B1I1 NETTRAN_DUMMY_6076 NETTRAN_DUMMY_6077 CLKBUF_X1 
XCLKBUF_X1_G2B1I33 n76 n76_G2B1I3 NETTRAN_DUMMY_6078 NETTRAN_DUMMY_6079 CLKBUF_X1 
XCLKBUF_X1_G2B1I43 n76 n76_G2B1I4 NETTRAN_DUMMY_6080 NETTRAN_DUMMY_6081 CLKBUF_X1 
XCLKBUF_X1_G2B1I24 clk_G1B1I2 n82_G2B1I2 NETTRAN_DUMMY_6082 NETTRAN_DUMMY_6083 CLKBUF_X1 
XCLKBUF_X1_G2B1I34 clk_G1B1I2 n82_G2B1I3 NETTRAN_DUMMY_6084 NETTRAN_DUMMY_6085 CLKBUF_X1 
XCLKBUF_X1_G2B1I44 clk_G1B1I2 n82_G2B1I4 NETTRAN_DUMMY_6086 NETTRAN_DUMMY_6087 CLKBUF_X1 
XCLKBUF_X1_G2B1I53 clk_G1B1I2 n82_G2B1I5 NETTRAN_DUMMY_6088 NETTRAN_DUMMY_6089 CLKBUF_X1 
XCLKBUF_X1_G2B1I63 clk_G1B1I2 n82_G2B1I6 NETTRAN_DUMMY_6090 NETTRAN_DUMMY_6091 CLKBUF_X1 
XCLKBUF_X1_G2B1I71 clk_G1B1I2 n82_G2B1I7 NETTRAN_DUMMY_6092 NETTRAN_DUMMY_6093 CLKBUF_X1 
XCLKBUF_X1_G2B1I81 clk_G1B1I2 n82_G2B1I8 NETTRAN_DUMMY_6094 NETTRAN_DUMMY_6095 CLKBUF_X1 
XCLKBUF_X1_G2B1I15 n80 n80_G2B1I1 NETTRAN_DUMMY_6096 NETTRAN_DUMMY_6097 CLKBUF_X1 
XCLKBUF_X1_G2B1I25 n80 n80_G2B1I2 NETTRAN_DUMMY_6098 NETTRAN_DUMMY_6099 CLKBUF_X1 
XCLKBUF_X1_G2B1I45 n80 n80_G2B1I4 NETTRAN_DUMMY_6100 NETTRAN_DUMMY_6101 CLKBUF_X1 
XCLKBUF_X1_G2B1I54 n80 n80_G2B1I5 NETTRAN_DUMMY_6102 NETTRAN_DUMMY_6103 CLKBUF_X1 
XCLKBUF_X1_G2B1I64 n80 n80_G2B1I6 NETTRAN_DUMMY_6104 NETTRAN_DUMMY_6105 CLKBUF_X1 
XCLKBUF_X1_G2B1I72 n80 n80_G2B1I7 NETTRAN_DUMMY_6106 NETTRAN_DUMMY_6107 CLKBUF_X1 
XU6 clk_cts_3 n125 NETTRAN_DUMMY_6108 NETTRAN_DUMMY_6109 CLKBUF_X1 
XCLKBUF_X3_G1B1I6 clk clk_G1B1I6 NETTRAN_DUMMY_6110 NETTRAN_DUMMY_6111 CLKBUF_X1 
XCLKBUF_X3_G1B1I3 clk clk_G1B1I3 NETTRAN_DUMMY_6112 NETTRAN_DUMMY_6113 CLKBUF_X1 
XU1 clk_G1B1I3 n76 NETTRAN_DUMMY_6114 NETTRAN_DUMMY_6115 CLKBUF_X1 
XCLKBUF_X2_G1B1I2 clk clk_G1B1I2 NETTRAN_DUMMY_6116 NETTRAN_DUMMY_6117 CLKBUF_X1 
XU5 clk_G1B1I3 n84 NETTRAN_DUMMY_6118 NETTRAN_DUMMY_6119 CLKBUF_X1 
XU2 clk_G1B1I6 n78 NETTRAN_DUMMY_6120 NETTRAN_DUMMY_6121 CLKBUF_X1 
XU3 clk_G1B1I6 n80 NETTRAN_DUMMY_6122 NETTRAN_DUMMY_6123 CLKBUF_X1 
XU4 n810 n304 NETTRAN_DUMMY_6124 NETTRAN_DUMMY_6125 BUF_X1 
XU8 n841 n305 NETTRAN_DUMMY_6126 NETTRAN_DUMMY_6127 BUF_X1 
XU23 n876 n306 NETTRAN_DUMMY_6128 NETTRAN_DUMMY_6129 BUF_X1 
XU24 n572 n307 NETTRAN_DUMMY_6130 NETTRAN_DUMMY_6131 BUF_X1 
XU25 n991 n308 NETTRAN_DUMMY_6132 NETTRAN_DUMMY_6133 BUF_X1 
XU26 n574 n309 NETTRAN_DUMMY_6134 NETTRAN_DUMMY_6135 BUF_X1 
XU27 n1018 n552 NETTRAN_DUMMY_6136 NETTRAN_DUMMY_6137 BUF_X1 
XU28 n1107 n553 NETTRAN_DUMMY_6138 NETTRAN_DUMMY_6139 BUF_X1 
XU29 n575 n554 NETTRAN_DUMMY_6140 NETTRAN_DUMMY_6141 BUF_X1 
XU30 n1150 n555 NETTRAN_DUMMY_6142 NETTRAN_DUMMY_6143 BUF_X1 
XU223 n1901 n556 NETTRAN_DUMMY_6144 NETTRAN_DUMMY_6145 BUF_X1 
XU468 n61 n1973 NETTRAN_DUMMY_6146 NETTRAN_DUMMY_6147 INV_X16 
XU469 n148 n1572 NETTRAN_DUMMY_6148 NETTRAN_DUMMY_6149 INV_X16 
XU470 n343 n1108 NETTRAN_DUMMY_6150 NETTRAN_DUMMY_6151 BUF_X1 
XU471 n3050 n1012 NETTRAN_DUMMY_6152 NETTRAN_DUMMY_6153 BUF_X1 
XU472 n990 n991 NETTRAN_DUMMY_6154 NETTRAN_DUMMY_6155 INV_X8 
XU473 n961 n962 NETTRAN_DUMMY_6156 NETTRAN_DUMMY_6157 INV_X8 
XU474 n911 n912 NETTRAN_DUMMY_6158 NETTRAN_DUMMY_6159 INV_X2 
XU475 n753 n557 NETTRAN_DUMMY_6160 NETTRAN_DUMMY_6161 INV_X1 
XU476 n557 n558 NETTRAN_DUMMY_6162 NETTRAN_DUMMY_6163 INV_X8 
XU477 n758 n559 NETTRAN_DUMMY_6164 NETTRAN_DUMMY_6165 BUF_X1 
XU478 n763 n560 NETTRAN_DUMMY_6166 NETTRAN_DUMMY_6167 CLKBUF_X1 
XU479 n773 n561 NETTRAN_DUMMY_6168 NETTRAN_DUMMY_6169 BUF_X1 
XU480 n772 n562 NETTRAN_DUMMY_6170 NETTRAN_DUMMY_6171 CLKBUF_X1 
XU481 n779 n563 NETTRAN_DUMMY_6172 NETTRAN_DUMMY_6173 BUF_X1 
XU482 n784 n564 NETTRAN_DUMMY_6174 NETTRAN_DUMMY_6175 BUF_X1 
XU483 n789 n565 NETTRAN_DUMMY_6176 NETTRAN_DUMMY_6177 BUF_X1 
XU484 n786 n566 NETTRAN_DUMMY_6178 NETTRAN_DUMMY_6179 CLKBUF_X1 
XU485 n794 n567 NETTRAN_DUMMY_6180 NETTRAN_DUMMY_6181 BUF_X1 
XU486 n791 n568 NETTRAN_DUMMY_6182 NETTRAN_DUMMY_6183 CLKBUF_X1 
XU487 n799 n569 NETTRAN_DUMMY_6184 NETTRAN_DUMMY_6185 INV_X1 
XU488 n569 n570 NETTRAN_DUMMY_6186 NETTRAN_DUMMY_6187 INV_X32 
XU489 n804 n571 NETTRAN_DUMMY_6188 NETTRAN_DUMMY_6189 BUF_X1 
XU490 n912 n572 NETTRAN_DUMMY_6190 NETTRAN_DUMMY_6191 BUF_X1 
XU491 n930 n573 NETTRAN_DUMMY_6192 NETTRAN_DUMMY_6193 BUF_X1 
XU492 n1014 n574 NETTRAN_DUMMY_6194 NETTRAN_DUMMY_6195 BUF_X1 
XU493 n1112 n575 NETTRAN_DUMMY_6196 NETTRAN_DUMMY_6197 BUF_X1 
XU494 z1_next[63] n576 NETTRAN_DUMMY_6198 NETTRAN_DUMMY_6199 CLKBUF_X1 
XU495 n1157 n577 NETTRAN_DUMMY_6200 NETTRAN_DUMMY_6201 BUF_X1 
XU496 n1162 n578 NETTRAN_DUMMY_6202 NETTRAN_DUMMY_6203 BUF_X1 
XU497 n1159 n579 NETTRAN_DUMMY_6204 NETTRAN_DUMMY_6205 CLKBUF_X1 
XU498 n1167 n580 NETTRAN_DUMMY_6206 NETTRAN_DUMMY_6207 INV_X1 
XU499 n580 n581 NETTRAN_DUMMY_6208 NETTRAN_DUMMY_6209 INV_X8 
XU500 n1178 n582 NETTRAN_DUMMY_6210 NETTRAN_DUMMY_6211 BUF_X1 
XU501 n1183 n583 NETTRAN_DUMMY_6212 NETTRAN_DUMMY_6213 BUF_X1 
XU502 n1188 n584 NETTRAN_DUMMY_6214 NETTRAN_DUMMY_6215 BUF_X1 
XU503 n1186 n585 NETTRAN_DUMMY_6216 NETTRAN_DUMMY_6217 CLKBUF_X1 
XU504 n1193 n586 NETTRAN_DUMMY_6218 NETTRAN_DUMMY_6219 BUF_X1 
XU505 n108 n587 NETTRAN_DUMMY_6220 NETTRAN_DUMMY_6221 CLKBUF_X1 
XU506 n1198 n588 NETTRAN_DUMMY_6222 NETTRAN_DUMMY_6223 CLKBUF_X1 
XU507 n1203 n589 NETTRAN_DUMMY_6224 NETTRAN_DUMMY_6225 BUF_X1 
XU508 n1208 n590 NETTRAN_DUMMY_6226 NETTRAN_DUMMY_6227 BUF_X1 
XU509 n1213 n591 NETTRAN_DUMMY_6228 NETTRAN_DUMMY_6229 BUF_X1 
XU510 n1218 n592 NETTRAN_DUMMY_6230 NETTRAN_DUMMY_6231 INV_X1 
XU511 n592 n593 NETTRAN_DUMMY_6232 NETTRAN_DUMMY_6233 INV_X8 
XU512 n1223 n594 NETTRAN_DUMMY_6234 NETTRAN_DUMMY_6235 BUF_X1 
XU513 n1220 n595 NETTRAN_DUMMY_6236 NETTRAN_DUMMY_6237 CLKBUF_X1 
XU514 n1233 n596 NETTRAN_DUMMY_6238 NETTRAN_DUMMY_6239 BUF_X1 
XU515 n114 n597 NETTRAN_DUMMY_6240 NETTRAN_DUMMY_6241 CLKBUF_X1 
XU516 n1243 n598 NETTRAN_DUMMY_6242 NETTRAN_DUMMY_6243 BUF_X1 
XU517 n1248 n599 NETTRAN_DUMMY_6244 NETTRAN_DUMMY_6245 BUF_X1 
XU518 n1246 n600 NETTRAN_DUMMY_6246 NETTRAN_DUMMY_6247 CLKBUF_X1 
XU519 n1259 n601 NETTRAN_DUMMY_6248 NETTRAN_DUMMY_6249 BUF_X1 
XU520 n1270 n602 NETTRAN_DUMMY_6250 NETTRAN_DUMMY_6251 BUF_X1 
XU521 n1268 n603 NETTRAN_DUMMY_6252 NETTRAN_DUMMY_6253 CLKBUF_X1 
XU522 n1275 n604 NETTRAN_DUMMY_6254 NETTRAN_DUMMY_6255 BUF_X1 
XU523 n1280 n605 NETTRAN_DUMMY_6256 NETTRAN_DUMMY_6257 BUF_X1 
XU524 n1285 n606 NETTRAN_DUMMY_6258 NETTRAN_DUMMY_6259 BUF_X1 
XU525 n1290 n607 NETTRAN_DUMMY_6260 NETTRAN_DUMMY_6261 CLKBUF_X1 
XU526 n1299 n608 NETTRAN_DUMMY_6262 NETTRAN_DUMMY_6263 BUF_X1 
XU527 n116 n609 NETTRAN_DUMMY_6264 NETTRAN_DUMMY_6265 CLKBUF_X1 
XU528 n1298 n610 NETTRAN_DUMMY_6266 NETTRAN_DUMMY_6267 CLKBUF_X1 
XU529 n1305 n611 NETTRAN_DUMMY_6268 NETTRAN_DUMMY_6269 BUF_X1 
XU530 n1310 n612 NETTRAN_DUMMY_6270 NETTRAN_DUMMY_6271 INV_X1 
XU531 n612 n613 NETTRAN_DUMMY_6272 NETTRAN_DUMMY_6273 INV_X8 
XU532 n1315 n614 NETTRAN_DUMMY_6274 NETTRAN_DUMMY_6275 BUF_X1 
XU533 n1320 n615 NETTRAN_DUMMY_6276 NETTRAN_DUMMY_6277 CLKBUF_X1 
XU534 n1325 n616 NETTRAN_DUMMY_6278 NETTRAN_DUMMY_6279 BUF_X1 
XU535 n1330 n617 NETTRAN_DUMMY_6280 NETTRAN_DUMMY_6281 BUF_X1 
XU536 n1328 n618 NETTRAN_DUMMY_6282 NETTRAN_DUMMY_6283 CLKBUF_X1 
XU537 n1335 n627 NETTRAN_DUMMY_6284 NETTRAN_DUMMY_6285 BUF_X1 
XU538 n1340 n628 NETTRAN_DUMMY_6286 NETTRAN_DUMMY_6287 BUF_X1 
XU539 n1345 n629 NETTRAN_DUMMY_6288 NETTRAN_DUMMY_6289 BUF_X1 
XU540 n1350 n630 NETTRAN_DUMMY_6290 NETTRAN_DUMMY_6291 BUF_X1 
XU541 n1347 n631 NETTRAN_DUMMY_6292 NETTRAN_DUMMY_6293 CLKBUF_X1 
XU542 n1355 n632 NETTRAN_DUMMY_6294 NETTRAN_DUMMY_6295 BUF_X1 
XU543 n1360 n633 NETTRAN_DUMMY_6296 NETTRAN_DUMMY_6297 CLKBUF_X1 
XU544 n1365 n634 NETTRAN_DUMMY_6298 NETTRAN_DUMMY_6299 BUF_X1 
XU545 n1370 n635 NETTRAN_DUMMY_6300 NETTRAN_DUMMY_6301 CLKBUF_X1 
XU546 n1373 n636 NETTRAN_DUMMY_6302 NETTRAN_DUMMY_6303 BUF_X1 
XU547 n1375 n637 NETTRAN_DUMMY_6304 NETTRAN_DUMMY_6305 CLKBUF_X1 
XU548 n1380 n638 NETTRAN_DUMMY_6306 NETTRAN_DUMMY_6307 BUF_X1 
XU549 n1385 n639 NETTRAN_DUMMY_6308 NETTRAN_DUMMY_6309 BUF_X1 
XU550 n1395 n640 NETTRAN_DUMMY_6310 NETTRAN_DUMMY_6311 INV_X1 
XU551 n640 n641 NETTRAN_DUMMY_6312 NETTRAN_DUMMY_6313 INV_X32 
XU552 n1405 n642 NETTRAN_DUMMY_6314 NETTRAN_DUMMY_6315 BUF_X1 
XU553 n158 n643 NETTRAN_DUMMY_6316 NETTRAN_DUMMY_6317 BUF_X1 
XU554 n1404 n644 NETTRAN_DUMMY_6318 NETTRAN_DUMMY_6319 CLKBUF_X1 
XU555 n1411 n645 NETTRAN_DUMMY_6320 NETTRAN_DUMMY_6321 BUF_X1 
XU556 n1427 n646 NETTRAN_DUMMY_6322 NETTRAN_DUMMY_6323 BUF_X1 
XU557 n1432 n647 NETTRAN_DUMMY_6324 NETTRAN_DUMMY_6325 BUF_X1 
XU558 n1437 n648 NETTRAN_DUMMY_6326 NETTRAN_DUMMY_6327 BUF_X1 
XU559 n1448 n649 NETTRAN_DUMMY_6328 NETTRAN_DUMMY_6329 BUF_X1 
XU560 n1459 n650 NETTRAN_DUMMY_6330 NETTRAN_DUMMY_6331 BUF_X1 
XU561 n1469 n651 NETTRAN_DUMMY_6332 NETTRAN_DUMMY_6333 BUF_X1 
XU562 n1468 n652 NETTRAN_DUMMY_6334 NETTRAN_DUMMY_6335 CLKBUF_X1 
XU563 n1475 n653 NETTRAN_DUMMY_6336 NETTRAN_DUMMY_6337 BUF_X1 
XU564 n1480 n654 NETTRAN_DUMMY_6338 NETTRAN_DUMMY_6339 BUF_X1 
XU565 n1488 n655 NETTRAN_DUMMY_6340 NETTRAN_DUMMY_6341 INV_X1 
XU566 n655 n656 NETTRAN_DUMMY_6342 NETTRAN_DUMMY_6343 INV_X32 
XU567 n1496 n657 NETTRAN_DUMMY_6344 NETTRAN_DUMMY_6345 BUF_X1 
XU568 n1501 n658 NETTRAN_DUMMY_6346 NETTRAN_DUMMY_6347 BUF_X1 
XU569 n1506 n659 NETTRAN_DUMMY_6348 NETTRAN_DUMMY_6349 BUF_X1 
XU570 n1511 n660 NETTRAN_DUMMY_6350 NETTRAN_DUMMY_6351 INV_X1 
XU571 n660 n661 NETTRAN_DUMMY_6352 NETTRAN_DUMMY_6353 INV_X8 
XU572 n1516 n662 NETTRAN_DUMMY_6354 NETTRAN_DUMMY_6355 BUF_X1 
XU573 n1521 n663 NETTRAN_DUMMY_6356 NETTRAN_DUMMY_6357 BUF_X1 
XU574 n1526 n664 NETTRAN_DUMMY_6358 NETTRAN_DUMMY_6359 INV_X1 
XU575 n664 n665 NETTRAN_DUMMY_6360 NETTRAN_DUMMY_6361 INV_X16 
XU576 n1531 n666 NETTRAN_DUMMY_6362 NETTRAN_DUMMY_6363 BUF_X1 
XU577 n181 n667 NETTRAN_DUMMY_6364 NETTRAN_DUMMY_6365 CLKBUF_X1 
XU578 n1542 n668 NETTRAN_DUMMY_6366 NETTRAN_DUMMY_6367 BUF_X1 
XU579 n1547 n669 NETTRAN_DUMMY_6368 NETTRAN_DUMMY_6369 BUF_X1 
XU580 n1552 n670 NETTRAN_DUMMY_6370 NETTRAN_DUMMY_6371 INV_X1 
XU581 n670 n671 NETTRAN_DUMMY_6372 NETTRAN_DUMMY_6373 INV_X8 
XU582 n1575 n672 NETTRAN_DUMMY_6374 NETTRAN_DUMMY_6375 BUF_X1 
XU583 n1574 n673 NETTRAN_DUMMY_6376 NETTRAN_DUMMY_6377 CLKBUF_X1 
XU584 n1592 n674 NETTRAN_DUMMY_6378 NETTRAN_DUMMY_6379 BUF_X1 
XU585 n1597 n675 NETTRAN_DUMMY_6380 NETTRAN_DUMMY_6381 BUF_X1 
XU586 n1602 n676 NETTRAN_DUMMY_6382 NETTRAN_DUMMY_6383 INV_X1 
XU587 n676 n677 NETTRAN_DUMMY_6384 NETTRAN_DUMMY_6385 INV_X8 
XU588 n1611 n678 NETTRAN_DUMMY_6386 NETTRAN_DUMMY_6387 BUF_X1 
XU589 n1618 n679 NETTRAN_DUMMY_6388 NETTRAN_DUMMY_6389 BUF_X1 
XU590 n1623 n680 NETTRAN_DUMMY_6390 NETTRAN_DUMMY_6391 BUF_X1 
XU591 n1639 n681 NETTRAN_DUMMY_6392 NETTRAN_DUMMY_6393 BUF_X1 
XU592 n1638 n682 NETTRAN_DUMMY_6394 NETTRAN_DUMMY_6395 CLKBUF_X1 
XU593 n1651 n683 NETTRAN_DUMMY_6396 NETTRAN_DUMMY_6397 BUF_X1 
XU594 n1656 n684 NETTRAN_DUMMY_6398 NETTRAN_DUMMY_6399 BUF_X1 
XU595 n1661 n685 NETTRAN_DUMMY_6400 NETTRAN_DUMMY_6401 BUF_X1 
XU596 n1666 n686 NETTRAN_DUMMY_6402 NETTRAN_DUMMY_6403 BUF_X1 
XU597 n1671 n687 NETTRAN_DUMMY_6404 NETTRAN_DUMMY_6405 BUF_X1 
XU598 n1675 n688 NETTRAN_DUMMY_6406 NETTRAN_DUMMY_6407 BUF_X1 
XU599 n1674 n689 NETTRAN_DUMMY_6408 NETTRAN_DUMMY_6409 CLKBUF_X1 
XU600 n1678 n690 NETTRAN_DUMMY_6410 NETTRAN_DUMMY_6411 BUF_X1 
XU601 n1677 n691 NETTRAN_DUMMY_6412 NETTRAN_DUMMY_6413 CLKBUF_X1 
XU602 n1686 n692 NETTRAN_DUMMY_6414 NETTRAN_DUMMY_6415 BUF_X1 
XU603 n1697 n693 NETTRAN_DUMMY_6416 NETTRAN_DUMMY_6417 BUF_X1 
XU604 n1702 n694 NETTRAN_DUMMY_6418 NETTRAN_DUMMY_6419 BUF_X1 
XU605 n1713 n695 NETTRAN_DUMMY_6420 NETTRAN_DUMMY_6421 BUF_X1 
XU606 n1716 n696 NETTRAN_DUMMY_6422 NETTRAN_DUMMY_6423 CLKBUF_X1 
XU607 n1728 n697 NETTRAN_DUMMY_6424 NETTRAN_DUMMY_6425 BUF_X1 
XU608 n54 n698 NETTRAN_DUMMY_6426 NETTRAN_DUMMY_6427 CLKBUF_X1 
XU609 n1727 n699 NETTRAN_DUMMY_6428 NETTRAN_DUMMY_6429 CLKBUF_X1 
XU610 n33 n700 NETTRAN_DUMMY_6430 NETTRAN_DUMMY_6431 BUF_X1 
XU611 n26 n701 NETTRAN_DUMMY_6432 NETTRAN_DUMMY_6433 BUF_X1 
XU612 n1755 n702 NETTRAN_DUMMY_6434 NETTRAN_DUMMY_6435 BUF_X1 
XU613 n19 n703 NETTRAN_DUMMY_6436 NETTRAN_DUMMY_6437 BUF_X1 
XU614 n1760 n704 NETTRAN_DUMMY_6438 NETTRAN_DUMMY_6439 CLKBUF_X1 
XU615 n1762 n705 NETTRAN_DUMMY_6440 NETTRAN_DUMMY_6441 BUF_X1 
XU616 n1761 n706 NETTRAN_DUMMY_6442 NETTRAN_DUMMY_6443 CLKBUF_X1 
XU617 n1770 n707 NETTRAN_DUMMY_6444 NETTRAN_DUMMY_6445 BUF_X1 
XU618 n1781 n708 NETTRAN_DUMMY_6446 NETTRAN_DUMMY_6447 BUF_X1 
XU619 n1786 n709 NETTRAN_DUMMY_6448 NETTRAN_DUMMY_6449 BUF_X1 
XU620 n1795 n710 NETTRAN_DUMMY_6450 NETTRAN_DUMMY_6451 BUF_X1 
XU621 n1802 n711 NETTRAN_DUMMY_6452 NETTRAN_DUMMY_6453 CLKBUF_X1 
XU622 n1813 n712 NETTRAN_DUMMY_6454 NETTRAN_DUMMY_6455 BUF_X1 
XU623 n1818 n713 NETTRAN_DUMMY_6456 NETTRAN_DUMMY_6457 BUF_X1 
XU624 n1823 n714 NETTRAN_DUMMY_6458 NETTRAN_DUMMY_6459 BUF_X1 
XU625 n1828 n715 NETTRAN_DUMMY_6460 NETTRAN_DUMMY_6461 BUF_X1 
XU626 n1833 n716 NETTRAN_DUMMY_6462 NETTRAN_DUMMY_6463 BUF_X1 
XU627 n1844 n717 NETTRAN_DUMMY_6464 NETTRAN_DUMMY_6465 CLKBUF_X1 
XU628 n1852 n718 NETTRAN_DUMMY_6466 NETTRAN_DUMMY_6467 BUF_X1 
XU629 n49 n719 NETTRAN_DUMMY_6468 NETTRAN_DUMMY_6469 CLKBUF_X1 
XU630 n1859 n720 NETTRAN_DUMMY_6470 NETTRAN_DUMMY_6471 BUF_X1 
XU631 n1868 n721 NETTRAN_DUMMY_6472 NETTRAN_DUMMY_6473 BUF_X1 
XU632 n1875 n722 NETTRAN_DUMMY_6474 NETTRAN_DUMMY_6475 BUF_X1 
XU633 n1878 n723 NETTRAN_DUMMY_6476 NETTRAN_DUMMY_6477 CLKBUF_X1 
XU634 n1885 n724 NETTRAN_DUMMY_6478 NETTRAN_DUMMY_6479 BUF_X1 
XU635 n1884 n725 NETTRAN_DUMMY_6480 NETTRAN_DUMMY_6481 CLKBUF_X1 
XU636 n45 n726 NETTRAN_DUMMY_6482 NETTRAN_DUMMY_6483 BUF_X1 
XU637 n38 n727 NETTRAN_DUMMY_6484 NETTRAN_DUMMY_6485 BUF_X1 
XU638 n1904 n728 NETTRAN_DUMMY_6486 NETTRAN_DUMMY_6487 BUF_X1 
XU639 n31 n729 NETTRAN_DUMMY_6488 NETTRAN_DUMMY_6489 BUF_X1 
XU640 n1911 n730 NETTRAN_DUMMY_6490 NETTRAN_DUMMY_6491 BUF_X1 
XU641 n1916 n731 NETTRAN_DUMMY_6492 NETTRAN_DUMMY_6493 BUF_X1 
XU642 n17 n732 NETTRAN_DUMMY_6494 NETTRAN_DUMMY_6495 BUF_X1 
XU643 n1921 n733 NETTRAN_DUMMY_6496 NETTRAN_DUMMY_6497 CLKBUF_X1 
XU644 n1930 n734 NETTRAN_DUMMY_6498 NETTRAN_DUMMY_6499 BUF_X1 
XU645 n123 n735 NETTRAN_DUMMY_6500 NETTRAN_DUMMY_6501 CLKBUF_X1 
XU646 n1929 n736 NETTRAN_DUMMY_6502 NETTRAN_DUMMY_6503 CLKBUF_X1 
XU647 n1942 n737 NETTRAN_DUMMY_6504 NETTRAN_DUMMY_6505 INV_X1 
XU648 n737 n738 NETTRAN_DUMMY_6506 NETTRAN_DUMMY_6507 INV_X4 
XU649 n1947 n739 NETTRAN_DUMMY_6508 NETTRAN_DUMMY_6509 BUF_X1 
XU650 n1958 n740 NETTRAN_DUMMY_6510 NETTRAN_DUMMY_6511 BUF_X1 
XU651 n1963 n741 NETTRAN_DUMMY_6512 NETTRAN_DUMMY_6513 BUF_X1 
XU652 n1968 n742 NETTRAN_DUMMY_6514 NETTRAN_DUMMY_6515 CLKBUF_X1 
XU653 n1972 n743 NETTRAN_DUMMY_6516 NETTRAN_DUMMY_6517 INV_X1 
XU654 n743 n744 NETTRAN_DUMMY_6518 NETTRAN_DUMMY_6519 INV_X32 
XU655 n1985 n745 NETTRAN_DUMMY_6520 NETTRAN_DUMMY_6521 BUF_X1 
XU656 n1990 n746 NETTRAN_DUMMY_6522 NETTRAN_DUMMY_6523 BUF_X1 
XU657 n1995 n747 NETTRAN_DUMMY_6524 NETTRAN_DUMMY_6525 BUF_X1 
XU658 n2012 n748 NETTRAN_DUMMY_6526 NETTRAN_DUMMY_6527 BUF_X1 
XU659 n752 n749 NETTRAN_DUMMY_6528 NETTRAN_DUMMY_6529 CLKBUF_X1 
XU660 n749 n750 NETTRAN_DUMMY_6530 NETTRAN_DUMMY_6531 INV_X32 
XU661 n750 n751 NETTRAN_DUMMY_6532 NETTRAN_DUMMY_6533 INV_X1 
XU662 n402 n752 NETTRAN_DUMMY_6534 NETTRAN_DUMMY_6535 INV_X1 
XU663 n751 n753 NETTRAN_DUMMY_6536 NETTRAN_DUMMY_6537 INV_X32 
XU664 n757 n754 NETTRAN_DUMMY_6538 NETTRAN_DUMMY_6539 CLKBUF_X1 
XU665 n754 n755 NETTRAN_DUMMY_6540 NETTRAN_DUMMY_6541 INV_X32 
XU666 n755 n756 NETTRAN_DUMMY_6542 NETTRAN_DUMMY_6543 INV_X1 
XU667 n389 n757 NETTRAN_DUMMY_6544 NETTRAN_DUMMY_6545 INV_X1 
XU668 n756 n758 NETTRAN_DUMMY_6546 NETTRAN_DUMMY_6547 INV_X32 
XU669 n762 n759 NETTRAN_DUMMY_6548 NETTRAN_DUMMY_6549 CLKBUF_X1 
XU670 n759 n760 NETTRAN_DUMMY_6550 NETTRAN_DUMMY_6551 INV_X32 
XU671 n760 n761 NETTRAN_DUMMY_6552 NETTRAN_DUMMY_6553 INV_X1 
XU672 n376 n762 NETTRAN_DUMMY_6554 NETTRAN_DUMMY_6555 INV_X1 
XU673 n761 n763 NETTRAN_DUMMY_6556 NETTRAN_DUMMY_6557 INV_X32 
XU674 n769 n764 NETTRAN_DUMMY_6558 NETTRAN_DUMMY_6559 INV_X1 
XU675 n764 n765 NETTRAN_DUMMY_6560 NETTRAN_DUMMY_6561 INV_X32 
XU676 n768 n766 NETTRAN_DUMMY_6562 NETTRAN_DUMMY_6563 INV_X32 
XU677 n766 n767 NETTRAN_DUMMY_6564 NETTRAN_DUMMY_6565 INV_X1 
XU678 n421 n768 NETTRAN_DUMMY_6566 NETTRAN_DUMMY_6567 INV_X1 
XU679 n767 n769 NETTRAN_DUMMY_6568 NETTRAN_DUMMY_6569 INV_X32 
XU680 n408 n770 NETTRAN_DUMMY_6570 NETTRAN_DUMMY_6571 INV_X1 
XU681 n770 n771 NETTRAN_DUMMY_6572 NETTRAN_DUMMY_6573 INV_X32 
XU682 n771 n772 NETTRAN_DUMMY_6574 NETTRAN_DUMMY_6575 INV_X1 
XU683 n562 n773 NETTRAN_DUMMY_6576 NETTRAN_DUMMY_6577 INV_X32 
XU684 n159 n774 NETTRAN_DUMMY_6578 NETTRAN_DUMMY_6579 CLKBUF_X1 
XU685 n778 n775 NETTRAN_DUMMY_6580 NETTRAN_DUMMY_6581 CLKBUF_X1 
XU686 n775 n776 NETTRAN_DUMMY_6582 NETTRAN_DUMMY_6583 INV_X32 
XU687 n776 n777 NETTRAN_DUMMY_6584 NETTRAN_DUMMY_6585 INV_X1 
XU688 n395 n778 NETTRAN_DUMMY_6586 NETTRAN_DUMMY_6587 INV_X1 
XU689 n777 n779 NETTRAN_DUMMY_6588 NETTRAN_DUMMY_6589 INV_X32 
XU690 n783 n780 NETTRAN_DUMMY_6590 NETTRAN_DUMMY_6591 CLKBUF_X1 
XU691 n382 n781 NETTRAN_DUMMY_6592 NETTRAN_DUMMY_6593 INV_X1 
XU692 n781 n782 NETTRAN_DUMMY_6594 NETTRAN_DUMMY_6595 INV_X32 
XU693 n782 n783 NETTRAN_DUMMY_6596 NETTRAN_DUMMY_6597 INV_X1 
XU694 n780 n784 NETTRAN_DUMMY_6598 NETTRAN_DUMMY_6599 INV_X32 
XU695 n788 n785 NETTRAN_DUMMY_6600 NETTRAN_DUMMY_6601 CLKBUF_X1 
XU696 n785 n786 NETTRAN_DUMMY_6602 NETTRAN_DUMMY_6603 INV_X32 
XU697 n566 n787 NETTRAN_DUMMY_6604 NETTRAN_DUMMY_6605 INV_X1 
XU698 n427 n788 NETTRAN_DUMMY_6606 NETTRAN_DUMMY_6607 INV_X1 
XU699 n787 n789 NETTRAN_DUMMY_6608 NETTRAN_DUMMY_6609 INV_X32 
XU700 n793 n790 NETTRAN_DUMMY_6610 NETTRAN_DUMMY_6611 CLKBUF_X1 
XU701 n790 n791 NETTRAN_DUMMY_6612 NETTRAN_DUMMY_6613 INV_X32 
XU702 n568 n792 NETTRAN_DUMMY_6614 NETTRAN_DUMMY_6615 INV_X1 
XU703 n414 n793 NETTRAN_DUMMY_6616 NETTRAN_DUMMY_6617 INV_X1 
XU704 n792 n794 NETTRAN_DUMMY_6618 NETTRAN_DUMMY_6619 INV_X32 
XU705 n798 n795 NETTRAN_DUMMY_6620 NETTRAN_DUMMY_6621 CLKBUF_X1 
XU706 n795 n796 NETTRAN_DUMMY_6622 NETTRAN_DUMMY_6623 INV_X32 
XU707 n796 n797 NETTRAN_DUMMY_6624 NETTRAN_DUMMY_6625 INV_X1 
XU708 n401 n798 NETTRAN_DUMMY_6626 NETTRAN_DUMMY_6627 INV_X1 
XU709 n797 n799 NETTRAN_DUMMY_6628 NETTRAN_DUMMY_6629 INV_X32 
XU710 n803 n800 NETTRAN_DUMMY_6630 NETTRAN_DUMMY_6631 CLKBUF_X1 
XU711 n388 n801 NETTRAN_DUMMY_6632 NETTRAN_DUMMY_6633 INV_X1 
XU712 n801 n802 NETTRAN_DUMMY_6634 NETTRAN_DUMMY_6635 INV_X32 
XU713 n802 n803 NETTRAN_DUMMY_6636 NETTRAN_DUMMY_6637 INV_X1 
XU714 n800 n804 NETTRAN_DUMMY_6638 NETTRAN_DUMMY_6639 INV_X32 
XU715 n8 n805 NETTRAN_DUMMY_6640 NETTRAN_DUMMY_6641 INV_X1 
XU716 n805 n806 NETTRAN_DUMMY_6642 NETTRAN_DUMMY_6643 INV_X32 
XU717 n233 n807 NETTRAN_DUMMY_6644 NETTRAN_DUMMY_6645 INV_X1 
XU718 n807 n808 NETTRAN_DUMMY_6646 NETTRAN_DUMMY_6647 INV_X32 
XU719 N3091 n809 NETTRAN_DUMMY_6648 NETTRAN_DUMMY_6649 INV_X1 
XU720 n809 n810 NETTRAN_DUMMY_6650 NETTRAN_DUMMY_6651 INV_X32 
XU721 n816 n811 NETTRAN_DUMMY_6652 NETTRAN_DUMMY_6653 INV_X1 
XU723 n235 n813 NETTRAN_DUMMY_6654 NETTRAN_DUMMY_6655 INV_X1 
XU724 n813 n814 NETTRAN_DUMMY_6656 NETTRAN_DUMMY_6657 INV_X32 
XU725 N3081 n815 NETTRAN_DUMMY_6658 NETTRAN_DUMMY_6659 INV_X1 
XU726 n815 n816 NETTRAN_DUMMY_6660 NETTRAN_DUMMY_6661 INV_X32 
XU727 n822 n817 NETTRAN_DUMMY_6662 NETTRAN_DUMMY_6663 INV_X1 
XU728 n817 n818 NETTRAN_DUMMY_6664 NETTRAN_DUMMY_6665 INV_X16 
XU729 n237 n819 NETTRAN_DUMMY_6666 NETTRAN_DUMMY_6667 INV_X1 
XU730 n819 n820 NETTRAN_DUMMY_6668 NETTRAN_DUMMY_6669 INV_X32 
XU731 N3071 n821 NETTRAN_DUMMY_6670 NETTRAN_DUMMY_6671 INV_X1 
XU732 n821 n822 NETTRAN_DUMMY_6672 NETTRAN_DUMMY_6673 INV_X32 
XU733 n828 n823 NETTRAN_DUMMY_6674 NETTRAN_DUMMY_6675 INV_X1 
XU734 n823 n824 NETTRAN_DUMMY_6676 NETTRAN_DUMMY_6677 INV_X8 
XU735 n239 n825 NETTRAN_DUMMY_6678 NETTRAN_DUMMY_6679 INV_X1 
XU736 n825 n826 NETTRAN_DUMMY_6680 NETTRAN_DUMMY_6681 INV_X32 
XU737 N3061 n827 NETTRAN_DUMMY_6682 NETTRAN_DUMMY_6683 INV_X1 
XU738 n827 n828 NETTRAN_DUMMY_6684 NETTRAN_DUMMY_6685 INV_X32 
XU739 n834 n829 NETTRAN_DUMMY_6686 NETTRAN_DUMMY_6687 INV_X1 
XU740 n829 n830 NETTRAN_DUMMY_6688 NETTRAN_DUMMY_6689 INV_X8 
XU741 n241 n831 NETTRAN_DUMMY_6690 NETTRAN_DUMMY_6691 INV_X1 
XU742 n831 n832 NETTRAN_DUMMY_6692 NETTRAN_DUMMY_6693 INV_X32 
XU743 N3051 n833 NETTRAN_DUMMY_6694 NETTRAN_DUMMY_6695 INV_X1 
XU744 n833 n834 NETTRAN_DUMMY_6696 NETTRAN_DUMMY_6697 INV_X32 
XU745 n840 n835 NETTRAN_DUMMY_6698 NETTRAN_DUMMY_6699 INV_X1 
XU746 n835 n836 NETTRAN_DUMMY_6700 NETTRAN_DUMMY_6701 INV_X32 
XU747 n243 n837 NETTRAN_DUMMY_6702 NETTRAN_DUMMY_6703 INV_X1 
XU748 n837 n838 NETTRAN_DUMMY_6704 NETTRAN_DUMMY_6705 INV_X32 
XU749 N3041 n839 NETTRAN_DUMMY_6706 NETTRAN_DUMMY_6707 INV_X1 
XU750 n839 n840 NETTRAN_DUMMY_6708 NETTRAN_DUMMY_6709 INV_X32 
XU751 n845 n841 NETTRAN_DUMMY_6710 NETTRAN_DUMMY_6711 CLKBUF_X1 
XU752 n245 n842 NETTRAN_DUMMY_6712 NETTRAN_DUMMY_6713 INV_X1 
XU753 n842 n843 NETTRAN_DUMMY_6714 NETTRAN_DUMMY_6715 INV_X32 
XU754 N303 n844 NETTRAN_DUMMY_6716 NETTRAN_DUMMY_6717 INV_X1 
XU755 n844 n845 NETTRAN_DUMMY_6718 NETTRAN_DUMMY_6719 INV_X32 
XU756 n850 n846 NETTRAN_DUMMY_6720 NETTRAN_DUMMY_6721 BUF_X1 
XU757 n2470 n847 NETTRAN_DUMMY_6722 NETTRAN_DUMMY_6723 INV_X1 
XU758 n847 n848 NETTRAN_DUMMY_6724 NETTRAN_DUMMY_6725 INV_X32 
XU759 N302 n849 NETTRAN_DUMMY_6726 NETTRAN_DUMMY_6727 INV_X1 
XU760 n849 n850 NETTRAN_DUMMY_6728 NETTRAN_DUMMY_6729 INV_X32 
XU761 n856 n851 NETTRAN_DUMMY_6730 NETTRAN_DUMMY_6731 INV_X1 
XU762 n851 n852 NETTRAN_DUMMY_6732 NETTRAN_DUMMY_6733 INV_X32 
XU763 n2490 n853 NETTRAN_DUMMY_6734 NETTRAN_DUMMY_6735 INV_X1 
XU764 n853 n854 NETTRAN_DUMMY_6736 NETTRAN_DUMMY_6737 INV_X32 
XU765 N301 n855 NETTRAN_DUMMY_6738 NETTRAN_DUMMY_6739 INV_X1 
XU766 n855 n856 NETTRAN_DUMMY_6740 NETTRAN_DUMMY_6741 INV_X32 
XU767 n862 n857 NETTRAN_DUMMY_6742 NETTRAN_DUMMY_6743 INV_X1 
XU768 n857 n858 NETTRAN_DUMMY_6744 NETTRAN_DUMMY_6745 INV_X32 
XU769 n2510 n859 NETTRAN_DUMMY_6746 NETTRAN_DUMMY_6747 INV_X1 
XU770 n859 n860 NETTRAN_DUMMY_6748 NETTRAN_DUMMY_6749 INV_X32 
XU771 N300 n861 NETTRAN_DUMMY_6750 NETTRAN_DUMMY_6751 INV_X1 
XU772 n861 n862 NETTRAN_DUMMY_6752 NETTRAN_DUMMY_6753 INV_X32 
XU773 n866 n863 NETTRAN_DUMMY_6754 NETTRAN_DUMMY_6755 INV_X1 
XU774 n863 n864 NETTRAN_DUMMY_6756 NETTRAN_DUMMY_6757 INV_X16 
XU775 N299 n865 NETTRAN_DUMMY_6758 NETTRAN_DUMMY_6759 INV_X1 
XU776 n865 n866 NETTRAN_DUMMY_6760 NETTRAN_DUMMY_6761 INV_X32 
XU777 n2530 n867 NETTRAN_DUMMY_6762 NETTRAN_DUMMY_6763 INV_X1 
XU778 n867 n868 NETTRAN_DUMMY_6764 NETTRAN_DUMMY_6765 INV_X32 
XU779 n872 n869 NETTRAN_DUMMY_6766 NETTRAN_DUMMY_6767 INV_X1 
XU780 n869 n870 NETTRAN_DUMMY_6768 NETTRAN_DUMMY_6769 INV_X16 
XU781 N298 n871 NETTRAN_DUMMY_6770 NETTRAN_DUMMY_6771 INV_X1 
XU782 n871 n872 NETTRAN_DUMMY_6772 NETTRAN_DUMMY_6773 INV_X32 
XU783 n25500 n873 NETTRAN_DUMMY_6774 NETTRAN_DUMMY_6775 INV_X1 
XU784 n873 n874 NETTRAN_DUMMY_6776 NETTRAN_DUMMY_6777 INV_X32 
XU785 n880 n875 NETTRAN_DUMMY_6778 NETTRAN_DUMMY_6779 INV_X1 
XU786 n875 n876 NETTRAN_DUMMY_6780 NETTRAN_DUMMY_6781 INV_X8 
XU787 n25700 n877 NETTRAN_DUMMY_6782 NETTRAN_DUMMY_6783 INV_X1 
XU788 n877 n878 NETTRAN_DUMMY_6784 NETTRAN_DUMMY_6785 INV_X32 
XU789 N297 n879 NETTRAN_DUMMY_6786 NETTRAN_DUMMY_6787 INV_X1 
XU790 n879 n880 NETTRAN_DUMMY_6788 NETTRAN_DUMMY_6789 INV_X32 
XU791 n884 n881 NETTRAN_DUMMY_6790 NETTRAN_DUMMY_6791 INV_X1 
XU792 n881 n882 NETTRAN_DUMMY_6792 NETTRAN_DUMMY_6793 INV_X16 
XU793 N296 n883 NETTRAN_DUMMY_6794 NETTRAN_DUMMY_6795 INV_X1 
XU794 n883 n884 NETTRAN_DUMMY_6796 NETTRAN_DUMMY_6797 INV_X32 
XU795 n25900 n885 NETTRAN_DUMMY_6798 NETTRAN_DUMMY_6799 INV_X1 
XU796 n885 n886 NETTRAN_DUMMY_6800 NETTRAN_DUMMY_6801 INV_X32 
XU797 n892 n887 NETTRAN_DUMMY_6802 NETTRAN_DUMMY_6803 INV_X1 
XU798 n887 n888 NETTRAN_DUMMY_6804 NETTRAN_DUMMY_6805 INV_X8 
XU799 n26100 n889 NETTRAN_DUMMY_6806 NETTRAN_DUMMY_6807 INV_X1 
XU800 n889 n890 NETTRAN_DUMMY_6808 NETTRAN_DUMMY_6809 INV_X32 
XU801 N295 n891 NETTRAN_DUMMY_6810 NETTRAN_DUMMY_6811 INV_X1 
XU802 n891 n892 NETTRAN_DUMMY_6812 NETTRAN_DUMMY_6813 INV_X32 
XU803 n898 n893 NETTRAN_DUMMY_6814 NETTRAN_DUMMY_6815 INV_X1 
XU804 n893 n894 NETTRAN_DUMMY_6816 NETTRAN_DUMMY_6817 INV_X16 
XU805 n2630 n895 NETTRAN_DUMMY_6818 NETTRAN_DUMMY_6819 INV_X1 
XU806 n895 n896 NETTRAN_DUMMY_6820 NETTRAN_DUMMY_6821 INV_X32 
XU807 N294 n897 NETTRAN_DUMMY_6822 NETTRAN_DUMMY_6823 INV_X1 
XU808 n897 n898 NETTRAN_DUMMY_6824 NETTRAN_DUMMY_6825 INV_X32 
XU809 n904 n899 NETTRAN_DUMMY_6826 NETTRAN_DUMMY_6827 INV_X1 
XU810 n899 n900 NETTRAN_DUMMY_6828 NETTRAN_DUMMY_6829 INV_X8 
XU811 n2650 n901 NETTRAN_DUMMY_6830 NETTRAN_DUMMY_6831 INV_X1 
XU812 n901 n902 NETTRAN_DUMMY_6832 NETTRAN_DUMMY_6833 INV_X32 
XU813 N293 n903 NETTRAN_DUMMY_6834 NETTRAN_DUMMY_6835 INV_X1 
XU814 n903 n904 NETTRAN_DUMMY_6836 NETTRAN_DUMMY_6837 INV_X32 
XU815 n910 n905 NETTRAN_DUMMY_6838 NETTRAN_DUMMY_6839 INV_X1 
XU816 n905 n906 NETTRAN_DUMMY_6840 NETTRAN_DUMMY_6841 INV_X16 
XU817 n2670 n907 NETTRAN_DUMMY_6842 NETTRAN_DUMMY_6843 INV_X1 
XU818 n907 n908 NETTRAN_DUMMY_6844 NETTRAN_DUMMY_6845 INV_X32 
XU819 N292 n909 NETTRAN_DUMMY_6846 NETTRAN_DUMMY_6847 INV_X1 
XU820 n909 n910 NETTRAN_DUMMY_6848 NETTRAN_DUMMY_6849 INV_X32 
XU821 n916 n911 NETTRAN_DUMMY_6850 NETTRAN_DUMMY_6851 INV_X1 
XU822 n2690 n913 NETTRAN_DUMMY_6852 NETTRAN_DUMMY_6853 INV_X1 
XU823 n913 n914 NETTRAN_DUMMY_6854 NETTRAN_DUMMY_6855 INV_X32 
XU824 N291 n915 NETTRAN_DUMMY_6856 NETTRAN_DUMMY_6857 INV_X1 
XU825 n915 n916 NETTRAN_DUMMY_6858 NETTRAN_DUMMY_6859 INV_X32 
XU826 n922 n917 NETTRAN_DUMMY_6860 NETTRAN_DUMMY_6861 INV_X1 
XU827 n917 n918 NETTRAN_DUMMY_6862 NETTRAN_DUMMY_6863 INV_X8 
XU828 n2710 n919 NETTRAN_DUMMY_6864 NETTRAN_DUMMY_6865 INV_X1 
XU829 n919 n920 NETTRAN_DUMMY_6866 NETTRAN_DUMMY_6867 INV_X32 
XU830 N290 n921 NETTRAN_DUMMY_6868 NETTRAN_DUMMY_6869 INV_X1 
XU831 n921 n922 NETTRAN_DUMMY_6870 NETTRAN_DUMMY_6871 INV_X32 
XU832 n928 n923 NETTRAN_DUMMY_6872 NETTRAN_DUMMY_6873 INV_X1 
XU833 n923 n924 NETTRAN_DUMMY_6874 NETTRAN_DUMMY_6875 INV_X16 
XU834 n2730 n925 NETTRAN_DUMMY_6876 NETTRAN_DUMMY_6877 INV_X1 
XU835 n925 n926 NETTRAN_DUMMY_6878 NETTRAN_DUMMY_6879 INV_X32 
XU836 N289 n927 NETTRAN_DUMMY_6880 NETTRAN_DUMMY_6881 INV_X1 
XU837 n927 n928 NETTRAN_DUMMY_6882 NETTRAN_DUMMY_6883 INV_X32 
XU838 n934 n929 NETTRAN_DUMMY_6884 NETTRAN_DUMMY_6885 INV_X1 
XU839 n929 n930 NETTRAN_DUMMY_6886 NETTRAN_DUMMY_6887 INV_X32 
XU840 n2750 n931 NETTRAN_DUMMY_6888 NETTRAN_DUMMY_6889 INV_X1 
XU841 n931 n932 NETTRAN_DUMMY_6890 NETTRAN_DUMMY_6891 INV_X32 
XU842 N288 n933 NETTRAN_DUMMY_6892 NETTRAN_DUMMY_6893 INV_X1 
XU843 n933 n934 NETTRAN_DUMMY_6894 NETTRAN_DUMMY_6895 INV_X32 
XU844 N287 n935 NETTRAN_DUMMY_6896 NETTRAN_DUMMY_6897 INV_X1 
XU845 n935 n936 NETTRAN_DUMMY_6898 NETTRAN_DUMMY_6899 INV_X32 
XU846 n2770 n937 NETTRAN_DUMMY_6900 NETTRAN_DUMMY_6901 INV_X1 
XU847 n937 n938 NETTRAN_DUMMY_6902 NETTRAN_DUMMY_6903 INV_X32 
XU848 n2790 n939 NETTRAN_DUMMY_6904 NETTRAN_DUMMY_6905 INV_X1 
XU849 n939 n940 NETTRAN_DUMMY_6906 NETTRAN_DUMMY_6907 INV_X32 
XU850 N286 n941 NETTRAN_DUMMY_6908 NETTRAN_DUMMY_6909 INV_X1 
XU851 n941 n942 NETTRAN_DUMMY_6910 NETTRAN_DUMMY_6911 INV_X32 
XU852 n948 n943 NETTRAN_DUMMY_6912 NETTRAN_DUMMY_6913 INV_X1 
XU853 n943 n944 NETTRAN_DUMMY_6914 NETTRAN_DUMMY_6915 INV_X16 
XU854 n2810 n945 NETTRAN_DUMMY_6916 NETTRAN_DUMMY_6917 INV_X1 
XU855 n945 n946 NETTRAN_DUMMY_6918 NETTRAN_DUMMY_6919 INV_X32 
XU856 N285 n947 NETTRAN_DUMMY_6920 NETTRAN_DUMMY_6921 INV_X1 
XU857 n947 n948 NETTRAN_DUMMY_6922 NETTRAN_DUMMY_6923 INV_X32 
XU858 n954 n949 NETTRAN_DUMMY_6924 NETTRAN_DUMMY_6925 INV_X1 
XU859 n949 n950 NETTRAN_DUMMY_6926 NETTRAN_DUMMY_6927 INV_X16 
XU860 n2830 n951 NETTRAN_DUMMY_6928 NETTRAN_DUMMY_6929 INV_X1 
XU861 n951 n952 NETTRAN_DUMMY_6930 NETTRAN_DUMMY_6931 INV_X32 
XU862 N284 n953 NETTRAN_DUMMY_6932 NETTRAN_DUMMY_6933 INV_X1 
XU863 n953 n954 NETTRAN_DUMMY_6934 NETTRAN_DUMMY_6935 INV_X32 
XU864 n960 n955 NETTRAN_DUMMY_6936 NETTRAN_DUMMY_6937 INV_X1 
XU865 n955 n956 NETTRAN_DUMMY_6938 NETTRAN_DUMMY_6939 INV_X8 
XU866 n2850 n957 NETTRAN_DUMMY_6940 NETTRAN_DUMMY_6941 INV_X1 
XU867 n957 n958 NETTRAN_DUMMY_6942 NETTRAN_DUMMY_6943 INV_X32 
XU868 N283 n959 NETTRAN_DUMMY_6944 NETTRAN_DUMMY_6945 INV_X1 
XU869 n959 n960 NETTRAN_DUMMY_6946 NETTRAN_DUMMY_6947 INV_X32 
XU870 n966 n961 NETTRAN_DUMMY_6948 NETTRAN_DUMMY_6949 INV_X1 
XU871 n2870 n963 NETTRAN_DUMMY_6950 NETTRAN_DUMMY_6951 INV_X1 
XU872 n963 n964 NETTRAN_DUMMY_6952 NETTRAN_DUMMY_6953 INV_X32 
XU873 N282 n965 NETTRAN_DUMMY_6954 NETTRAN_DUMMY_6955 INV_X1 
XU874 n965 n966 NETTRAN_DUMMY_6956 NETTRAN_DUMMY_6957 INV_X32 
XU875 n972 n967 NETTRAN_DUMMY_6958 NETTRAN_DUMMY_6959 INV_X1 
XU876 n967 n968 NETTRAN_DUMMY_6960 NETTRAN_DUMMY_6961 INV_X32 
XU877 n2890 n969 NETTRAN_DUMMY_6962 NETTRAN_DUMMY_6963 INV_X1 
XU878 n969 n970 NETTRAN_DUMMY_6964 NETTRAN_DUMMY_6965 INV_X32 
XU879 N281 n971 NETTRAN_DUMMY_6966 NETTRAN_DUMMY_6967 INV_X1 
XU880 n971 n972 NETTRAN_DUMMY_6968 NETTRAN_DUMMY_6969 INV_X32 
XU881 n975 n973 NETTRAN_DUMMY_6970 NETTRAN_DUMMY_6971 BUF_X1 
XU882 N280 n974 NETTRAN_DUMMY_6972 NETTRAN_DUMMY_6973 INV_X1 
XU883 n974 n975 NETTRAN_DUMMY_6974 NETTRAN_DUMMY_6975 INV_X32 
XU884 n2910 n976 NETTRAN_DUMMY_6976 NETTRAN_DUMMY_6977 INV_X1 
XU885 n976 n977 NETTRAN_DUMMY_6978 NETTRAN_DUMMY_6979 INV_X32 
XU886 n983 n978 NETTRAN_DUMMY_6980 NETTRAN_DUMMY_6981 INV_X1 
XU887 n978 n979 NETTRAN_DUMMY_6982 NETTRAN_DUMMY_6983 INV_X16 
XU888 n2930 n980 NETTRAN_DUMMY_6984 NETTRAN_DUMMY_6985 INV_X1 
XU889 n980 n981 NETTRAN_DUMMY_6986 NETTRAN_DUMMY_6987 INV_X32 
XU890 N279 n982 NETTRAN_DUMMY_6988 NETTRAN_DUMMY_6989 INV_X1 
XU891 n982 n983 NETTRAN_DUMMY_6990 NETTRAN_DUMMY_6991 INV_X32 
XU892 n989 n984 NETTRAN_DUMMY_6992 NETTRAN_DUMMY_6993 INV_X1 
XU893 n984 n985 NETTRAN_DUMMY_6994 NETTRAN_DUMMY_6995 INV_X16 
XU894 n2950 n986 NETTRAN_DUMMY_6996 NETTRAN_DUMMY_6997 INV_X1 
XU895 n986 n987 NETTRAN_DUMMY_6998 NETTRAN_DUMMY_6999 INV_X32 
XU896 N278 n988 NETTRAN_DUMMY_7000 NETTRAN_DUMMY_7001 INV_X1 
XU897 n988 n989 NETTRAN_DUMMY_7002 NETTRAN_DUMMY_7003 INV_X32 
XU898 n995 n990 NETTRAN_DUMMY_7004 NETTRAN_DUMMY_7005 INV_X1 
XU899 n2970 n992 NETTRAN_DUMMY_7006 NETTRAN_DUMMY_7007 INV_X1 
XU900 n992 n993 NETTRAN_DUMMY_7008 NETTRAN_DUMMY_7009 INV_X32 
XU901 N277 n994 NETTRAN_DUMMY_7010 NETTRAN_DUMMY_7011 INV_X1 
XU902 n994 n995 NETTRAN_DUMMY_7012 NETTRAN_DUMMY_7013 INV_X32 
XU903 n1001 n996 NETTRAN_DUMMY_7014 NETTRAN_DUMMY_7015 INV_X1 
XU904 n996 n997 NETTRAN_DUMMY_7016 NETTRAN_DUMMY_7017 INV_X16 
XU905 n2990 n998 NETTRAN_DUMMY_7018 NETTRAN_DUMMY_7019 INV_X1 
XU906 n998 n999 NETTRAN_DUMMY_7020 NETTRAN_DUMMY_7021 INV_X32 
XU907 N276 n1000 NETTRAN_DUMMY_7022 NETTRAN_DUMMY_7023 INV_X1 
XU908 n1000 n1001 NETTRAN_DUMMY_7024 NETTRAN_DUMMY_7025 INV_X32 
XU909 n1005 n1002 NETTRAN_DUMMY_7026 NETTRAN_DUMMY_7027 INV_X1 
XU910 n1002 n1003 NETTRAN_DUMMY_7028 NETTRAN_DUMMY_7029 INV_X16 
XU911 N275 n1004 NETTRAN_DUMMY_7030 NETTRAN_DUMMY_7031 INV_X1 
XU912 n1004 n1005 NETTRAN_DUMMY_7032 NETTRAN_DUMMY_7033 INV_X32 
XU913 n3010 n1006 NETTRAN_DUMMY_7034 NETTRAN_DUMMY_7035 INV_X1 
XU914 n1006 n1007 NETTRAN_DUMMY_7036 NETTRAN_DUMMY_7037 INV_X32 
XU915 N274 n1008 NETTRAN_DUMMY_7038 NETTRAN_DUMMY_7039 INV_X1 
XU916 n1008 n1009 NETTRAN_DUMMY_7040 NETTRAN_DUMMY_7041 INV_X32 
XU917 n3030 n1010 NETTRAN_DUMMY_7042 NETTRAN_DUMMY_7043 INV_X1 
XU918 n1010 n1011 NETTRAN_DUMMY_7044 NETTRAN_DUMMY_7045 INV_X32 
XU919 N273 n1013 NETTRAN_DUMMY_7046 NETTRAN_DUMMY_7047 INV_X1 
XU920 n1013 n1014 NETTRAN_DUMMY_7048 NETTRAN_DUMMY_7049 INV_X32 
XU921 n1012 n1015 NETTRAN_DUMMY_7050 NETTRAN_DUMMY_7051 INV_X1 
XU922 n1015 n1016 NETTRAN_DUMMY_7052 NETTRAN_DUMMY_7053 INV_X32 
XU923 n1022 n1017 NETTRAN_DUMMY_7054 NETTRAN_DUMMY_7055 INV_X1 
XU924 n1017 n1018 NETTRAN_DUMMY_7056 NETTRAN_DUMMY_7057 INV_X16 
XU925 n3070 n1019 NETTRAN_DUMMY_7058 NETTRAN_DUMMY_7059 INV_X1 
XU926 n1019 n1020 NETTRAN_DUMMY_7060 NETTRAN_DUMMY_7061 INV_X32 
XU927 N272 n1021 NETTRAN_DUMMY_7062 NETTRAN_DUMMY_7063 INV_X1 
XU928 n1021 n1022 NETTRAN_DUMMY_7064 NETTRAN_DUMMY_7065 INV_X32 
XU929 n1027 n1023 NETTRAN_DUMMY_7066 NETTRAN_DUMMY_7067 BUF_X1 
XU930 n3090 n1024 NETTRAN_DUMMY_7068 NETTRAN_DUMMY_7069 INV_X1 
XU931 n1024 n1025 NETTRAN_DUMMY_7070 NETTRAN_DUMMY_7071 INV_X32 
XU932 N271 n1026 NETTRAN_DUMMY_7072 NETTRAN_DUMMY_7073 INV_X1 
XU933 n1026 n1027 NETTRAN_DUMMY_7074 NETTRAN_DUMMY_7075 INV_X32 
XU934 n1033 n1028 NETTRAN_DUMMY_7076 NETTRAN_DUMMY_7077 INV_X1 
XU935 n1028 n1029 NETTRAN_DUMMY_7078 NETTRAN_DUMMY_7079 INV_X16 
XU936 n311 n1030 NETTRAN_DUMMY_7080 NETTRAN_DUMMY_7081 INV_X1 
XU937 n1030 n1031 NETTRAN_DUMMY_7082 NETTRAN_DUMMY_7083 INV_X32 
XU938 N270 n1032 NETTRAN_DUMMY_7084 NETTRAN_DUMMY_7085 INV_X1 
XU939 n1032 n1033 NETTRAN_DUMMY_7086 NETTRAN_DUMMY_7087 INV_X32 
XU940 n1039 n1034 NETTRAN_DUMMY_7088 NETTRAN_DUMMY_7089 INV_X1 
XU941 n1034 n1035 NETTRAN_DUMMY_7090 NETTRAN_DUMMY_7091 INV_X32 
XU942 n313 n1036 NETTRAN_DUMMY_7092 NETTRAN_DUMMY_7093 INV_X1 
XU943 n1036 n1037 NETTRAN_DUMMY_7094 NETTRAN_DUMMY_7095 INV_X32 
XU944 N269 n1038 NETTRAN_DUMMY_7096 NETTRAN_DUMMY_7097 INV_X1 
XU945 n1038 n1039 NETTRAN_DUMMY_7098 NETTRAN_DUMMY_7099 INV_X32 
XU946 n1041 n1040 NETTRAN_DUMMY_7100 NETTRAN_DUMMY_7101 CLKBUF_X1 
XU947 n315 n1041 NETTRAN_DUMMY_7102 NETTRAN_DUMMY_7103 INV_X1 
XU948 n1040 n1042 NETTRAN_DUMMY_7104 NETTRAN_DUMMY_7105 INV_X32 
XU949 N268 n1043 NETTRAN_DUMMY_7106 NETTRAN_DUMMY_7107 INV_X1 
XU950 n1043 n1044 NETTRAN_DUMMY_7108 NETTRAN_DUMMY_7109 INV_X32 
XU951 n1049 n1045 NETTRAN_DUMMY_7110 NETTRAN_DUMMY_7111 BUF_X1 
XU952 n317 n1046 NETTRAN_DUMMY_7112 NETTRAN_DUMMY_7113 INV_X1 
XU953 n1046 n1047 NETTRAN_DUMMY_7114 NETTRAN_DUMMY_7115 INV_X32 
XU954 N267 n1048 NETTRAN_DUMMY_7116 NETTRAN_DUMMY_7117 INV_X1 
XU955 n1048 n1049 NETTRAN_DUMMY_7118 NETTRAN_DUMMY_7119 INV_X32 
XU956 n1055 n1050 NETTRAN_DUMMY_7120 NETTRAN_DUMMY_7121 INV_X1 
XU957 n1050 n1051 NETTRAN_DUMMY_7122 NETTRAN_DUMMY_7123 INV_X16 
XU958 n319 n1052 NETTRAN_DUMMY_7124 NETTRAN_DUMMY_7125 INV_X1 
XU959 n1052 n1053 NETTRAN_DUMMY_7126 NETTRAN_DUMMY_7127 INV_X32 
XU960 N266 n1054 NETTRAN_DUMMY_7128 NETTRAN_DUMMY_7129 INV_X1 
XU961 n1054 n1055 NETTRAN_DUMMY_7130 NETTRAN_DUMMY_7131 INV_X32 
XU962 n1060 n1056 NETTRAN_DUMMY_7132 NETTRAN_DUMMY_7133 BUF_X1 
XU963 n321 n1057 NETTRAN_DUMMY_7134 NETTRAN_DUMMY_7135 INV_X1 
XU964 n1057 n1058 NETTRAN_DUMMY_7136 NETTRAN_DUMMY_7137 INV_X32 
XU965 N265 n1059 NETTRAN_DUMMY_7138 NETTRAN_DUMMY_7139 INV_X1 
XU966 n1059 n1060 NETTRAN_DUMMY_7140 NETTRAN_DUMMY_7141 INV_X32 
XU967 n1062 n1061 NETTRAN_DUMMY_7142 NETTRAN_DUMMY_7143 CLKBUF_X1 
XU968 n323 n1062 NETTRAN_DUMMY_7144 NETTRAN_DUMMY_7145 INV_X1 
XU969 n1061 n1063 NETTRAN_DUMMY_7146 NETTRAN_DUMMY_7147 INV_X32 
XU970 N264 n1064 NETTRAN_DUMMY_7148 NETTRAN_DUMMY_7149 INV_X1 
XU971 n1064 n1065 NETTRAN_DUMMY_7150 NETTRAN_DUMMY_7151 INV_X32 
XU972 n1070 n1066 NETTRAN_DUMMY_7152 NETTRAN_DUMMY_7153 BUF_X1 
XU973 n325 n1067 NETTRAN_DUMMY_7154 NETTRAN_DUMMY_7155 INV_X1 
XU974 n1067 n1068 NETTRAN_DUMMY_7156 NETTRAN_DUMMY_7157 INV_X32 
XU975 N263 n1069 NETTRAN_DUMMY_7158 NETTRAN_DUMMY_7159 INV_X1 
XU976 n1069 n1070 NETTRAN_DUMMY_7160 NETTRAN_DUMMY_7161 INV_X32 
XU977 n1075 n1071 NETTRAN_DUMMY_7162 NETTRAN_DUMMY_7163 BUF_X1 
XU978 n327 n1072 NETTRAN_DUMMY_7164 NETTRAN_DUMMY_7165 INV_X1 
XU979 n1072 n1073 NETTRAN_DUMMY_7166 NETTRAN_DUMMY_7167 INV_X32 
XU980 N262 n1074 NETTRAN_DUMMY_7168 NETTRAN_DUMMY_7169 INV_X1 
XU981 n1074 n1075 NETTRAN_DUMMY_7170 NETTRAN_DUMMY_7171 INV_X32 
XU982 n1078 n1076 NETTRAN_DUMMY_7172 NETTRAN_DUMMY_7173 BUF_X1 
XU983 N2610 n1077 NETTRAN_DUMMY_7174 NETTRAN_DUMMY_7175 INV_X1 
XU984 n1077 n1078 NETTRAN_DUMMY_7176 NETTRAN_DUMMY_7177 INV_X32 
XU985 n329 n1079 NETTRAN_DUMMY_7178 NETTRAN_DUMMY_7179 INV_X1 
XU986 n1079 n1080 NETTRAN_DUMMY_7180 NETTRAN_DUMMY_7181 INV_X32 
XU987 n1084 n1081 NETTRAN_DUMMY_7182 NETTRAN_DUMMY_7183 INV_X1 
XU988 n1081 n1082 NETTRAN_DUMMY_7184 NETTRAN_DUMMY_7185 INV_X32 
XU989 N2600 n1083 NETTRAN_DUMMY_7186 NETTRAN_DUMMY_7187 INV_X1 
XU990 n1083 n1084 NETTRAN_DUMMY_7188 NETTRAN_DUMMY_7189 INV_X32 
XU991 n1088 n1085 NETTRAN_DUMMY_7190 NETTRAN_DUMMY_7191 INV_X1 
XU992 n1085 n1086 NETTRAN_DUMMY_7192 NETTRAN_DUMMY_7193 INV_X32 
XU993 N2590 n1087 NETTRAN_DUMMY_7194 NETTRAN_DUMMY_7195 INV_X1 
XU994 n1087 n1088 NETTRAN_DUMMY_7196 NETTRAN_DUMMY_7197 INV_X32 
XU995 n335 n1089 NETTRAN_DUMMY_7198 NETTRAN_DUMMY_7199 INV_X1 
XU996 n1089 n1090 NETTRAN_DUMMY_7200 NETTRAN_DUMMY_7201 INV_X32 
XU997 N2580 n1091 NETTRAN_DUMMY_7202 NETTRAN_DUMMY_7203 INV_X1 
XU998 n1091 n1092 NETTRAN_DUMMY_7204 NETTRAN_DUMMY_7205 INV_X32 
XU999 n1097 n1093 NETTRAN_DUMMY_7206 NETTRAN_DUMMY_7207 BUF_X1 
XU1000 n337 n1094 NETTRAN_DUMMY_7208 NETTRAN_DUMMY_7209 INV_X1 
XU1001 n1094 n1095 NETTRAN_DUMMY_7210 NETTRAN_DUMMY_7211 INV_X32 
XU1002 N2570 n1096 NETTRAN_DUMMY_7212 NETTRAN_DUMMY_7213 INV_X1 
XU1003 n1096 n1097 NETTRAN_DUMMY_7214 NETTRAN_DUMMY_7215 INV_X32 
XU1004 n1102 n1098 NETTRAN_DUMMY_7216 NETTRAN_DUMMY_7217 BUF_X1 
XU1005 n339 n1099 NETTRAN_DUMMY_7218 NETTRAN_DUMMY_7219 INV_X1 
XU1006 n1099 n1100 NETTRAN_DUMMY_7220 NETTRAN_DUMMY_7221 INV_X32 
XU1007 N2560 n1101 NETTRAN_DUMMY_7222 NETTRAN_DUMMY_7223 INV_X1 
XU1008 n1101 n1102 NETTRAN_DUMMY_7224 NETTRAN_DUMMY_7225 INV_X32 
XU1009 n1104 n1103 NETTRAN_DUMMY_7226 NETTRAN_DUMMY_7227 CLKBUF_X1 
XU1010 n341 n1104 NETTRAN_DUMMY_7228 NETTRAN_DUMMY_7229 INV_X1 
XU1011 n1103 n1105 NETTRAN_DUMMY_7230 NETTRAN_DUMMY_7231 INV_X32 
XU1012 N2550 n1106 NETTRAN_DUMMY_7232 NETTRAN_DUMMY_7233 INV_X1 
XU1013 n1106 n1107 NETTRAN_DUMMY_7234 NETTRAN_DUMMY_7235 INV_X32 
XU1014 n1108 n1109 NETTRAN_DUMMY_7236 NETTRAN_DUMMY_7237 INV_X1 
XU1015 n1109 n1110 NETTRAN_DUMMY_7238 NETTRAN_DUMMY_7239 INV_X32 
XU1016 N2540 n1111 NETTRAN_DUMMY_7240 NETTRAN_DUMMY_7241 INV_X1 
XU1017 n1111 n1112 NETTRAN_DUMMY_7242 NETTRAN_DUMMY_7243 INV_X32 
XU1018 n1114 n1113 NETTRAN_DUMMY_7244 NETTRAN_DUMMY_7245 CLKBUF_X1 
XU1019 n346 n1114 NETTRAN_DUMMY_7246 NETTRAN_DUMMY_7247 INV_X1 
XU1020 n1113 n1115 NETTRAN_DUMMY_7248 NETTRAN_DUMMY_7249 INV_X32 
XU1021 N253 n1116 NETTRAN_DUMMY_7250 NETTRAN_DUMMY_7251 INV_X1 
XU1022 n1116 n1117 NETTRAN_DUMMY_7252 NETTRAN_DUMMY_7253 INV_X32 
XU1023 n1122 n1118 NETTRAN_DUMMY_7254 NETTRAN_DUMMY_7255 BUF_X1 
XU1024 n349 n1119 NETTRAN_DUMMY_7256 NETTRAN_DUMMY_7257 INV_X1 
XU1025 n1119 n1120 NETTRAN_DUMMY_7258 NETTRAN_DUMMY_7259 INV_X32 
XU1026 N2520 n1121 NETTRAN_DUMMY_7260 NETTRAN_DUMMY_7261 INV_X1 
XU1027 n1121 n1122 NETTRAN_DUMMY_7262 NETTRAN_DUMMY_7263 INV_X32 
XU1028 n352 n1123 NETTRAN_DUMMY_7264 NETTRAN_DUMMY_7265 INV_X1 
XU1029 n1123 n1124 NETTRAN_DUMMY_7266 NETTRAN_DUMMY_7267 INV_X32 
XU1030 N251 n1125 NETTRAN_DUMMY_7268 NETTRAN_DUMMY_7269 INV_X1 
XU1031 n1125 n1126 NETTRAN_DUMMY_7270 NETTRAN_DUMMY_7271 INV_X32 
XU1032 n1131 n1127 NETTRAN_DUMMY_7272 NETTRAN_DUMMY_7273 BUF_X1 
XU1033 n356 n1128 NETTRAN_DUMMY_7274 NETTRAN_DUMMY_7275 INV_X1 
XU1034 n1128 n1129 NETTRAN_DUMMY_7276 NETTRAN_DUMMY_7277 INV_X32 
XU1035 N2500 n1130 NETTRAN_DUMMY_7278 NETTRAN_DUMMY_7279 INV_X1 
XU1036 n1130 n1131 NETTRAN_DUMMY_7280 NETTRAN_DUMMY_7281 INV_X32 
XU1037 n1136 n1132 NETTRAN_DUMMY_7282 NETTRAN_DUMMY_7283 BUF_X1 
XU1038 n360 n1133 NETTRAN_DUMMY_7284 NETTRAN_DUMMY_7285 INV_X1 
XU1039 n1133 n1134 NETTRAN_DUMMY_7286 NETTRAN_DUMMY_7287 INV_X32 
XU1040 N249 n1135 NETTRAN_DUMMY_7288 NETTRAN_DUMMY_7289 INV_X1 
XU1041 n1135 n1136 NETTRAN_DUMMY_7290 NETTRAN_DUMMY_7291 INV_X32 
XU1042 n1141 n1137 NETTRAN_DUMMY_7292 NETTRAN_DUMMY_7293 BUF_X1 
XU1043 n364 n1138 NETTRAN_DUMMY_7294 NETTRAN_DUMMY_7295 INV_X1 
XU1044 n1138 n1139 NETTRAN_DUMMY_7296 NETTRAN_DUMMY_7297 INV_X32 
XU1045 N2480 n1140 NETTRAN_DUMMY_7298 NETTRAN_DUMMY_7299 INV_X1 
XU1046 n1140 n1141 NETTRAN_DUMMY_7300 NETTRAN_DUMMY_7301 INV_X32 
XU1047 n1146 n1142 NETTRAN_DUMMY_7302 NETTRAN_DUMMY_7303 BUF_X1 
XU1048 n368 n1143 NETTRAN_DUMMY_7304 NETTRAN_DUMMY_7305 INV_X1 
XU1049 n1143 n1144 NETTRAN_DUMMY_7306 NETTRAN_DUMMY_7307 INV_X32 
XU1050 N247 n1145 NETTRAN_DUMMY_7308 NETTRAN_DUMMY_7309 INV_X1 
XU1051 n1145 n1146 NETTRAN_DUMMY_7310 NETTRAN_DUMMY_7311 INV_X32 
XU1052 n372 n1147 NETTRAN_DUMMY_7312 NETTRAN_DUMMY_7313 INV_X1 
XU1053 n1147 n1148 NETTRAN_DUMMY_7314 NETTRAN_DUMMY_7315 INV_X32 
XU1054 N2460 n1149 NETTRAN_DUMMY_7316 NETTRAN_DUMMY_7317 INV_X1 
XU1055 n1149 n1150 NETTRAN_DUMMY_7318 NETTRAN_DUMMY_7319 INV_X32 
XU1056 n164 n1151 NETTRAN_DUMMY_7320 NETTRAN_DUMMY_7321 INV_X32 
XU1057 n1151 n1152 NETTRAN_DUMMY_7322 NETTRAN_DUMMY_7323 INV_X1 
XU1058 n1156 n1153 NETTRAN_DUMMY_7324 NETTRAN_DUMMY_7325 CLKBUF_X1 
XU1059 n1153 n1154 NETTRAN_DUMMY_7326 NETTRAN_DUMMY_7327 INV_X32 
XU1060 n1154 n1155 NETTRAN_DUMMY_7328 NETTRAN_DUMMY_7329 INV_X1 
XU1061 n470 n1156 NETTRAN_DUMMY_7330 NETTRAN_DUMMY_7331 INV_X1 
XU1062 n1155 n1157 NETTRAN_DUMMY_7332 NETTRAN_DUMMY_7333 INV_X32 
XU1063 n1161 n1158 NETTRAN_DUMMY_7334 NETTRAN_DUMMY_7335 CLKBUF_X1 
XU1064 n1158 n1159 NETTRAN_DUMMY_7336 NETTRAN_DUMMY_7337 INV_X32 
XU1065 n579 n1160 NETTRAN_DUMMY_7338 NETTRAN_DUMMY_7339 INV_X1 
XU1066 n446 n1161 NETTRAN_DUMMY_7340 NETTRAN_DUMMY_7341 INV_X1 
XU1067 n1160 n1162 NETTRAN_DUMMY_7342 NETTRAN_DUMMY_7343 INV_X32 
XU1068 n1164 n1163 NETTRAN_DUMMY_7344 NETTRAN_DUMMY_7345 CLKBUF_X1 
XU1069 n480 n1164 NETTRAN_DUMMY_7346 NETTRAN_DUMMY_7347 INV_X1 
XU1070 n1163 n1165 NETTRAN_DUMMY_7348 NETTRAN_DUMMY_7349 INV_X32 
XU1071 n1165 n1166 NETTRAN_DUMMY_7350 NETTRAN_DUMMY_7351 INV_X1 
XU1072 n1166 n1167 NETTRAN_DUMMY_7352 NETTRAN_DUMMY_7353 INV_X32 
XU1073 n1173 n1168 NETTRAN_DUMMY_7354 NETTRAN_DUMMY_7355 INV_X1 
XU1074 n1168 n1169 NETTRAN_DUMMY_7356 NETTRAN_DUMMY_7357 INV_X32 
XU1075 n1172 n1170 NETTRAN_DUMMY_7358 NETTRAN_DUMMY_7359 INV_X32 
XU1076 n1170 n1171 NETTRAN_DUMMY_7360 NETTRAN_DUMMY_7361 INV_X1 
XU1077 n456 n1172 NETTRAN_DUMMY_7362 NETTRAN_DUMMY_7363 INV_X1 
XU1078 n1171 n1173 NETTRAN_DUMMY_7364 NETTRAN_DUMMY_7365 INV_X32 
XU1079 n1177 n1174 NETTRAN_DUMMY_7366 NETTRAN_DUMMY_7367 CLKBUF_X1 
XU1080 n1174 n1175 NETTRAN_DUMMY_7368 NETTRAN_DUMMY_7369 INV_X32 
XU1081 n1175 n1176 NETTRAN_DUMMY_7370 NETTRAN_DUMMY_7371 INV_X1 
XU1082 n495 n1177 NETTRAN_DUMMY_7372 NETTRAN_DUMMY_7373 INV_X1 
XU1083 n1176 n1178 NETTRAN_DUMMY_7374 NETTRAN_DUMMY_7375 INV_X32 
XU1084 n1182 n1179 NETTRAN_DUMMY_7376 NETTRAN_DUMMY_7377 CLKBUF_X1 
XU1085 n1179 n1180 NETTRAN_DUMMY_7378 NETTRAN_DUMMY_7379 INV_X32 
XU1086 n1180 n1181 NETTRAN_DUMMY_7380 NETTRAN_DUMMY_7381 INV_X1 
XU1087 n471 n1182 NETTRAN_DUMMY_7382 NETTRAN_DUMMY_7383 INV_X1 
XU1088 n1181 n1183 NETTRAN_DUMMY_7384 NETTRAN_DUMMY_7385 INV_X32 
XU1089 n1187 n1184 NETTRAN_DUMMY_7386 NETTRAN_DUMMY_7387 CLKBUF_X1 
XU1090 n447 n1185 NETTRAN_DUMMY_7388 NETTRAN_DUMMY_7389 INV_X1 
XU1091 n1185 n1186 NETTRAN_DUMMY_7390 NETTRAN_DUMMY_7391 INV_X32 
XU1092 n585 n1187 NETTRAN_DUMMY_7392 NETTRAN_DUMMY_7393 INV_X1 
XU1093 n1184 n1188 NETTRAN_DUMMY_7394 NETTRAN_DUMMY_7395 INV_X32 
XU1094 n1190 n1189 NETTRAN_DUMMY_7396 NETTRAN_DUMMY_7397 CLKBUF_X1 
XU1095 n481 n1190 NETTRAN_DUMMY_7398 NETTRAN_DUMMY_7399 INV_X1 
XU1096 n1189 n1191 NETTRAN_DUMMY_7400 NETTRAN_DUMMY_7401 INV_X32 
XU1097 n1191 n1192 NETTRAN_DUMMY_7402 NETTRAN_DUMMY_7403 INV_X1 
XU1098 n1192 n1193 NETTRAN_DUMMY_7404 NETTRAN_DUMMY_7405 INV_X32 
XU1099 n1197 n1194 NETTRAN_DUMMY_7406 NETTRAN_DUMMY_7407 CLKBUF_X1 
XU1100 n457 n1195 NETTRAN_DUMMY_7408 NETTRAN_DUMMY_7409 INV_X1 
XU1101 n1195 n1196 NETTRAN_DUMMY_7410 NETTRAN_DUMMY_7411 INV_X32 
XU1102 n1196 n1197 NETTRAN_DUMMY_7412 NETTRAN_DUMMY_7413 INV_X1 
XU1103 n1194 n1198 NETTRAN_DUMMY_7414 NETTRAN_DUMMY_7415 INV_X32 
XU1104 n1202 n1199 NETTRAN_DUMMY_7416 NETTRAN_DUMMY_7417 CLKBUF_X1 
XU1105 n1199 n1200 NETTRAN_DUMMY_7418 NETTRAN_DUMMY_7419 INV_X32 
XU1106 n1200 n1201 NETTRAN_DUMMY_7420 NETTRAN_DUMMY_7421 INV_X1 
XU1107 n491 n1202 NETTRAN_DUMMY_7422 NETTRAN_DUMMY_7423 INV_X1 
XU1108 n1201 n1203 NETTRAN_DUMMY_7424 NETTRAN_DUMMY_7425 INV_X32 
XU1109 n1207 n1204 NETTRAN_DUMMY_7426 NETTRAN_DUMMY_7427 CLKBUF_X1 
XU1110 n1204 n1205 NETTRAN_DUMMY_7428 NETTRAN_DUMMY_7429 INV_X32 
XU1111 n1205 n1206 NETTRAN_DUMMY_7430 NETTRAN_DUMMY_7431 INV_X1 
XU1112 n467 n1207 NETTRAN_DUMMY_7432 NETTRAN_DUMMY_7433 INV_X1 
XU1113 n1206 n1208 NETTRAN_DUMMY_7434 NETTRAN_DUMMY_7435 INV_X32 
XU1114 n1212 n1209 NETTRAN_DUMMY_7436 NETTRAN_DUMMY_7437 CLKBUF_X1 
XU1115 n1209 n1210 NETTRAN_DUMMY_7438 NETTRAN_DUMMY_7439 INV_X32 
XU1116 n1210 n1211 NETTRAN_DUMMY_7440 NETTRAN_DUMMY_7441 INV_X1 
XU1117 n443 n1212 NETTRAN_DUMMY_7442 NETTRAN_DUMMY_7443 INV_X1 
XU1118 n1211 n1213 NETTRAN_DUMMY_7444 NETTRAN_DUMMY_7445 INV_X32 
XU1119 n1217 n1214 NETTRAN_DUMMY_7446 NETTRAN_DUMMY_7447 CLKBUF_X1 
XU1120 n1214 n1215 NETTRAN_DUMMY_7448 NETTRAN_DUMMY_7449 INV_X32 
XU1121 n1215 n1216 NETTRAN_DUMMY_7450 NETTRAN_DUMMY_7451 INV_X1 
XU1122 n477 n1217 NETTRAN_DUMMY_7452 NETTRAN_DUMMY_7453 INV_X1 
XU1123 n1216 n1218 NETTRAN_DUMMY_7454 NETTRAN_DUMMY_7455 INV_X32 
XU1124 n1222 n1219 NETTRAN_DUMMY_7456 NETTRAN_DUMMY_7457 CLKBUF_X1 
XU1125 n1219 n1220 NETTRAN_DUMMY_7458 NETTRAN_DUMMY_7459 INV_X32 
XU1126 n595 n1221 NETTRAN_DUMMY_7460 NETTRAN_DUMMY_7461 INV_X1 
XU1127 n453 n1222 NETTRAN_DUMMY_7462 NETTRAN_DUMMY_7463 INV_X1 
XU1128 n1221 n1223 NETTRAN_DUMMY_7464 NETTRAN_DUMMY_7465 INV_X32 
XU1129 n1225 n1224 NETTRAN_DUMMY_7466 NETTRAN_DUMMY_7467 CLKBUF_X1 
XU1130 n487 n1225 NETTRAN_DUMMY_7468 NETTRAN_DUMMY_7469 INV_X1 
XU1131 n1224 n1226 NETTRAN_DUMMY_7470 NETTRAN_DUMMY_7471 INV_X32 
XU1132 n1226 n1227 NETTRAN_DUMMY_7472 NETTRAN_DUMMY_7473 INV_X1 
XU1133 n1227 n1228 NETTRAN_DUMMY_7474 NETTRAN_DUMMY_7475 INV_X32 
XU1134 n1230 n1229 NETTRAN_DUMMY_7476 NETTRAN_DUMMY_7477 CLKBUF_X1 
XU1135 n463 n1230 NETTRAN_DUMMY_7478 NETTRAN_DUMMY_7479 INV_X1 
XU1136 n1229 n1231 NETTRAN_DUMMY_7480 NETTRAN_DUMMY_7481 INV_X32 
XU1137 n1231 n1232 NETTRAN_DUMMY_7482 NETTRAN_DUMMY_7483 INV_X1 
XU1138 n1232 n1233 NETTRAN_DUMMY_7484 NETTRAN_DUMMY_7485 INV_X32 
XU1139 n1238 n1234 NETTRAN_DUMMY_7486 NETTRAN_DUMMY_7487 BUF_X1 
XU1140 n1237 n1235 NETTRAN_DUMMY_7488 NETTRAN_DUMMY_7489 INV_X32 
XU1141 n1235 n1236 NETTRAN_DUMMY_7490 NETTRAN_DUMMY_7491 INV_X1 
XU1142 n439 n1237 NETTRAN_DUMMY_7492 NETTRAN_DUMMY_7493 INV_X1 
XU1143 n1236 n1238 NETTRAN_DUMMY_7494 NETTRAN_DUMMY_7495 INV_X32 
XU1144 n1242 n1239 NETTRAN_DUMMY_7496 NETTRAN_DUMMY_7497 CLKBUF_X1 
XU1145 n1239 n1240 NETTRAN_DUMMY_7498 NETTRAN_DUMMY_7499 INV_X32 
XU1146 n1240 n1241 NETTRAN_DUMMY_7500 NETTRAN_DUMMY_7501 INV_X1 
XU1147 n473 n1242 NETTRAN_DUMMY_7502 NETTRAN_DUMMY_7503 INV_X1 
XU1148 n1241 n1243 NETTRAN_DUMMY_7504 NETTRAN_DUMMY_7505 INV_X32 
XU1149 n1247 n1244 NETTRAN_DUMMY_7506 NETTRAN_DUMMY_7507 CLKBUF_X1 
XU1150 n449 n1245 NETTRAN_DUMMY_7508 NETTRAN_DUMMY_7509 INV_X1 
XU1151 n1245 n1246 NETTRAN_DUMMY_7510 NETTRAN_DUMMY_7511 INV_X32 
XU1152 n600 n1247 NETTRAN_DUMMY_7512 NETTRAN_DUMMY_7513 INV_X1 
XU1153 n1244 n1248 NETTRAN_DUMMY_7514 NETTRAN_DUMMY_7515 INV_X32 
XU1154 n1254 n1249 NETTRAN_DUMMY_7516 NETTRAN_DUMMY_7517 INV_X1 
XU1155 n1249 n1250 NETTRAN_DUMMY_7518 NETTRAN_DUMMY_7519 INV_X32 
XU1156 n488 n1251 NETTRAN_DUMMY_7520 NETTRAN_DUMMY_7521 INV_X1 
XU1157 n1251 n1252 NETTRAN_DUMMY_7522 NETTRAN_DUMMY_7523 INV_X32 
XU1158 n1252 n1253 NETTRAN_DUMMY_7524 NETTRAN_DUMMY_7525 INV_X1 
XU1159 n1253 n1254 NETTRAN_DUMMY_7526 NETTRAN_DUMMY_7527 INV_X32 
XU1160 n1258 n1255 NETTRAN_DUMMY_7528 NETTRAN_DUMMY_7529 CLKBUF_X1 
XU1161 n1255 n1256 NETTRAN_DUMMY_7530 NETTRAN_DUMMY_7531 INV_X32 
XU1162 n1256 n1257 NETTRAN_DUMMY_7532 NETTRAN_DUMMY_7533 INV_X1 
XU1163 n464 n1258 NETTRAN_DUMMY_7534 NETTRAN_DUMMY_7535 INV_X1 
XU1164 n1257 n1259 NETTRAN_DUMMY_7536 NETTRAN_DUMMY_7537 INV_X32 
XU1165 n1265 n1260 NETTRAN_DUMMY_7538 NETTRAN_DUMMY_7539 INV_X1 
XU1166 n1260 n1261 NETTRAN_DUMMY_7540 NETTRAN_DUMMY_7541 INV_X32 
XU1167 n440 n1262 NETTRAN_DUMMY_7542 NETTRAN_DUMMY_7543 INV_X1 
XU1168 n1262 n1263 NETTRAN_DUMMY_7544 NETTRAN_DUMMY_7545 INV_X32 
XU1169 n1263 n1264 NETTRAN_DUMMY_7546 NETTRAN_DUMMY_7547 INV_X1 
XU1170 n1264 n1265 NETTRAN_DUMMY_7548 NETTRAN_DUMMY_7549 INV_X32 
XU1171 n1269 n1266 NETTRAN_DUMMY_7550 NETTRAN_DUMMY_7551 CLKBUF_X1 
XU1172 n483 n1267 NETTRAN_DUMMY_7552 NETTRAN_DUMMY_7553 INV_X1 
XU1173 n1267 n1268 NETTRAN_DUMMY_7554 NETTRAN_DUMMY_7555 INV_X32 
XU1174 n603 n1269 NETTRAN_DUMMY_7556 NETTRAN_DUMMY_7557 INV_X1 
XU1175 n1266 n1270 NETTRAN_DUMMY_7558 NETTRAN_DUMMY_7559 INV_X32 
XU1176 n1272 n1271 NETTRAN_DUMMY_7560 NETTRAN_DUMMY_7561 CLKBUF_X1 
XU1177 n459 n1272 NETTRAN_DUMMY_7562 NETTRAN_DUMMY_7563 INV_X1 
XU1178 n1271 n1273 NETTRAN_DUMMY_7564 NETTRAN_DUMMY_7565 INV_X32 
XU1179 n1273 n1274 NETTRAN_DUMMY_7566 NETTRAN_DUMMY_7567 INV_X1 
XU1180 n1274 n1275 NETTRAN_DUMMY_7568 NETTRAN_DUMMY_7569 INV_X32 
XU1181 n1279 n1276 NETTRAN_DUMMY_7570 NETTRAN_DUMMY_7571 CLKBUF_X1 
XU1182 n1276 n1277 NETTRAN_DUMMY_7572 NETTRAN_DUMMY_7573 INV_X32 
XU1183 n1277 n1278 NETTRAN_DUMMY_7574 NETTRAN_DUMMY_7575 INV_X1 
XU1184 n435 n1279 NETTRAN_DUMMY_7576 NETTRAN_DUMMY_7577 INV_X1 
XU1185 n1278 n1280 NETTRAN_DUMMY_7578 NETTRAN_DUMMY_7579 INV_X32 
XU1186 n1282 n1281 NETTRAN_DUMMY_7580 NETTRAN_DUMMY_7581 CLKBUF_X1 
XU1187 n474 n1282 NETTRAN_DUMMY_7582 NETTRAN_DUMMY_7583 INV_X1 
XU1188 n1281 n1283 NETTRAN_DUMMY_7584 NETTRAN_DUMMY_7585 INV_X32 
XU1189 n1283 n1284 NETTRAN_DUMMY_7586 NETTRAN_DUMMY_7587 INV_X1 
XU1190 n1284 n1285 NETTRAN_DUMMY_7588 NETTRAN_DUMMY_7589 INV_X32 
XU1191 n1289 n1286 NETTRAN_DUMMY_7590 NETTRAN_DUMMY_7591 CLKBUF_X1 
XU1192 n450 n1287 NETTRAN_DUMMY_7592 NETTRAN_DUMMY_7593 INV_X1 
XU1193 n1287 n1288 NETTRAN_DUMMY_7594 NETTRAN_DUMMY_7595 INV_X32 
XU1194 n1288 n1289 NETTRAN_DUMMY_7596 NETTRAN_DUMMY_7597 INV_X1 
XU1195 n1286 n1290 NETTRAN_DUMMY_7598 NETTRAN_DUMMY_7599 INV_X32 
XU1196 n1294 n1291 NETTRAN_DUMMY_7600 NETTRAN_DUMMY_7601 CLKBUF_X1 
XU1197 n1291 n1292 NETTRAN_DUMMY_7602 NETTRAN_DUMMY_7603 INV_X32 
XU1198 n1292 n1293 NETTRAN_DUMMY_7604 NETTRAN_DUMMY_7605 INV_X1 
XU1199 n489 n1294 NETTRAN_DUMMY_7606 NETTRAN_DUMMY_7607 INV_X1 
XU1200 n1293 n1295 NETTRAN_DUMMY_7608 NETTRAN_DUMMY_7609 INV_X32 
XU1201 n610 n1296 NETTRAN_DUMMY_7610 NETTRAN_DUMMY_7611 INV_X32 
XU1202 n1296 n1297 NETTRAN_DUMMY_7612 NETTRAN_DUMMY_7613 INV_X1 
XU1203 n465 n1298 NETTRAN_DUMMY_7614 NETTRAN_DUMMY_7615 INV_X1 
XU1204 n1297 n1299 NETTRAN_DUMMY_7616 NETTRAN_DUMMY_7617 INV_X32 
XU1205 n92 n1300 NETTRAN_DUMMY_7618 NETTRAN_DUMMY_7619 BUF_X1 
XU1206 n1304 n1301 NETTRAN_DUMMY_7620 NETTRAN_DUMMY_7621 CLKBUF_X1 
XU1207 n441 n1302 NETTRAN_DUMMY_7622 NETTRAN_DUMMY_7623 INV_X1 
XU1208 n1302 n1303 NETTRAN_DUMMY_7624 NETTRAN_DUMMY_7625 INV_X32 
XU1209 n1303 n1304 NETTRAN_DUMMY_7626 NETTRAN_DUMMY_7627 INV_X1 
XU1210 n1301 n1305 NETTRAN_DUMMY_7628 NETTRAN_DUMMY_7629 INV_X32 
XU1211 n1308 n1306 NETTRAN_DUMMY_7630 NETTRAN_DUMMY_7631 CLKBUF_X1 
XU1212 n1309 n1307 NETTRAN_DUMMY_7632 NETTRAN_DUMMY_7633 INV_X32 
XU1213 n1307 n1308 NETTRAN_DUMMY_7634 NETTRAN_DUMMY_7635 INV_X1 
XU1214 n484 n1309 NETTRAN_DUMMY_7636 NETTRAN_DUMMY_7637 INV_X1 
XU1215 n1306 n1310 NETTRAN_DUMMY_7638 NETTRAN_DUMMY_7639 INV_X32 
XU1216 n1314 n1311 NETTRAN_DUMMY_7640 NETTRAN_DUMMY_7641 CLKBUF_X1 
XU1217 n1311 n1312 NETTRAN_DUMMY_7642 NETTRAN_DUMMY_7643 INV_X32 
XU1218 n1312 n1313 NETTRAN_DUMMY_7644 NETTRAN_DUMMY_7645 INV_X1 
XU1219 n460 n1314 NETTRAN_DUMMY_7646 NETTRAN_DUMMY_7647 INV_X1 
XU1220 n1313 n1315 NETTRAN_DUMMY_7648 NETTRAN_DUMMY_7649 INV_X32 
XU1221 n1319 n1316 NETTRAN_DUMMY_7650 NETTRAN_DUMMY_7651 CLKBUF_X1 
XU1222 n1316 n1317 NETTRAN_DUMMY_7652 NETTRAN_DUMMY_7653 INV_X32 
XU1223 n1317 n1318 NETTRAN_DUMMY_7654 NETTRAN_DUMMY_7655 INV_X1 
XU1224 n436 n1319 NETTRAN_DUMMY_7656 NETTRAN_DUMMY_7657 INV_X1 
XU1225 n1318 n1320 NETTRAN_DUMMY_7658 NETTRAN_DUMMY_7659 INV_X32 
XU1226 n1324 n1321 NETTRAN_DUMMY_7660 NETTRAN_DUMMY_7661 CLKBUF_X1 
XU1227 n475 n1322 NETTRAN_DUMMY_7662 NETTRAN_DUMMY_7663 INV_X1 
XU1228 n1322 n1323 NETTRAN_DUMMY_7664 NETTRAN_DUMMY_7665 INV_X32 
XU1229 n1323 n1324 NETTRAN_DUMMY_7666 NETTRAN_DUMMY_7667 INV_X1 
XU1230 n1321 n1325 NETTRAN_DUMMY_7668 NETTRAN_DUMMY_7669 INV_X32 
XU1231 n1329 n1326 NETTRAN_DUMMY_7670 NETTRAN_DUMMY_7671 CLKBUF_X1 
XU1232 n451 n1327 NETTRAN_DUMMY_7672 NETTRAN_DUMMY_7673 INV_X1 
XU1233 n1327 n1328 NETTRAN_DUMMY_7674 NETTRAN_DUMMY_7675 INV_X32 
XU1234 n618 n1329 NETTRAN_DUMMY_7676 NETTRAN_DUMMY_7677 INV_X1 
XU1235 n1326 n1330 NETTRAN_DUMMY_7678 NETTRAN_DUMMY_7679 INV_X32 
XU1236 n1334 n1331 NETTRAN_DUMMY_7680 NETTRAN_DUMMY_7681 CLKBUF_X1 
XU1237 n1331 n1332 NETTRAN_DUMMY_7682 NETTRAN_DUMMY_7683 INV_X32 
XU1238 n1332 n1333 NETTRAN_DUMMY_7684 NETTRAN_DUMMY_7685 INV_X1 
XU1239 n490 n1334 NETTRAN_DUMMY_7686 NETTRAN_DUMMY_7687 INV_X1 
XU1240 n1333 n1335 NETTRAN_DUMMY_7688 NETTRAN_DUMMY_7689 INV_X32 
XU1241 n1339 n1336 NETTRAN_DUMMY_7690 NETTRAN_DUMMY_7691 CLKBUF_X1 
XU1242 n1336 n1337 NETTRAN_DUMMY_7692 NETTRAN_DUMMY_7693 INV_X32 
XU1243 n1337 n1338 NETTRAN_DUMMY_7694 NETTRAN_DUMMY_7695 INV_X1 
XU1244 n466 n1339 NETTRAN_DUMMY_7696 NETTRAN_DUMMY_7697 INV_X1 
XU1245 n1338 n1340 NETTRAN_DUMMY_7698 NETTRAN_DUMMY_7699 INV_X32 
XU1246 n1344 n1341 NETTRAN_DUMMY_7700 NETTRAN_DUMMY_7701 CLKBUF_X1 
XU1247 n1341 n1342 NETTRAN_DUMMY_7702 NETTRAN_DUMMY_7703 INV_X32 
XU1248 n1342 n1343 NETTRAN_DUMMY_7704 NETTRAN_DUMMY_7705 INV_X1 
XU1249 n442 n1344 NETTRAN_DUMMY_7706 NETTRAN_DUMMY_7707 INV_X1 
XU1250 n1343 n1345 NETTRAN_DUMMY_7708 NETTRAN_DUMMY_7709 INV_X32 
XU1251 n1349 n1346 NETTRAN_DUMMY_7710 NETTRAN_DUMMY_7711 CLKBUF_X1 
XU1252 n1346 n1347 NETTRAN_DUMMY_7712 NETTRAN_DUMMY_7713 INV_X32 
XU1253 n631 n1348 NETTRAN_DUMMY_7714 NETTRAN_DUMMY_7715 INV_X1 
XU1254 n485 n1349 NETTRAN_DUMMY_7716 NETTRAN_DUMMY_7717 INV_X1 
XU1255 n1348 n1350 NETTRAN_DUMMY_7718 NETTRAN_DUMMY_7719 INV_X32 
XU1256 n1354 n1351 NETTRAN_DUMMY_7720 NETTRAN_DUMMY_7721 CLKBUF_X1 
XU1257 n461 n1352 NETTRAN_DUMMY_7722 NETTRAN_DUMMY_7723 INV_X1 
XU1258 n1352 n1353 NETTRAN_DUMMY_7724 NETTRAN_DUMMY_7725 INV_X32 
XU1259 n1353 n1354 NETTRAN_DUMMY_7726 NETTRAN_DUMMY_7727 INV_X1 
XU1260 n1351 n1355 NETTRAN_DUMMY_7728 NETTRAN_DUMMY_7729 INV_X32 
XU1261 n1359 n1356 NETTRAN_DUMMY_7730 NETTRAN_DUMMY_7731 CLKBUF_X1 
XU1262 n437 n1357 NETTRAN_DUMMY_7732 NETTRAN_DUMMY_7733 INV_X1 
XU1263 n1357 n1358 NETTRAN_DUMMY_7734 NETTRAN_DUMMY_7735 INV_X32 
XU1264 n1358 n1359 NETTRAN_DUMMY_7736 NETTRAN_DUMMY_7737 INV_X1 
XU1265 n1356 n1360 NETTRAN_DUMMY_7738 NETTRAN_DUMMY_7739 INV_X32 
XU1266 n1364 n1361 NETTRAN_DUMMY_7740 NETTRAN_DUMMY_7741 CLKBUF_X1 
XU1267 n476 n1362 NETTRAN_DUMMY_7742 NETTRAN_DUMMY_7743 INV_X1 
XU1268 n1362 n1363 NETTRAN_DUMMY_7744 NETTRAN_DUMMY_7745 INV_X32 
XU1269 n1363 n1364 NETTRAN_DUMMY_7746 NETTRAN_DUMMY_7747 INV_X1 
XU1270 n1361 n1365 NETTRAN_DUMMY_7748 NETTRAN_DUMMY_7749 INV_X32 
XU1271 n1367 n1366 NETTRAN_DUMMY_7750 NETTRAN_DUMMY_7751 CLKBUF_X1 
XU1272 n452 n1367 NETTRAN_DUMMY_7752 NETTRAN_DUMMY_7753 INV_X1 
XU1273 n1366 n1368 NETTRAN_DUMMY_7754 NETTRAN_DUMMY_7755 INV_X32 
XU1274 n1368 n1369 NETTRAN_DUMMY_7756 NETTRAN_DUMMY_7757 INV_X1 
XU1275 n1369 n1370 NETTRAN_DUMMY_7758 NETTRAN_DUMMY_7759 INV_X32 
XU1276 n1372 n1371 NETTRAN_DUMMY_7760 NETTRAN_DUMMY_7761 CLKBUF_X1 
XU1277 n637 n1372 NETTRAN_DUMMY_7762 NETTRAN_DUMMY_7763 INV_X1 
XU1278 n1371 n1373 NETTRAN_DUMMY_7764 NETTRAN_DUMMY_7765 INV_X32 
XU1279 n486 n1374 NETTRAN_DUMMY_7766 NETTRAN_DUMMY_7767 INV_X1 
XU1280 n1374 n1375 NETTRAN_DUMMY_7768 NETTRAN_DUMMY_7769 INV_X32 
XU1281 n1379 n1376 NETTRAN_DUMMY_7770 NETTRAN_DUMMY_7771 CLKBUF_X1 
XU1282 n462 n1377 NETTRAN_DUMMY_7772 NETTRAN_DUMMY_7773 INV_X1 
XU1283 n1377 n1378 NETTRAN_DUMMY_7774 NETTRAN_DUMMY_7775 INV_X32 
XU1284 n1378 n1379 NETTRAN_DUMMY_7776 NETTRAN_DUMMY_7777 INV_X1 
XU1285 n1376 n1380 NETTRAN_DUMMY_7778 NETTRAN_DUMMY_7779 INV_X32 
XU1286 n1383 n1381 NETTRAN_DUMMY_7780 NETTRAN_DUMMY_7781 CLKBUF_X1 
XU1287 n1384 n1382 NETTRAN_DUMMY_7782 NETTRAN_DUMMY_7783 INV_X32 
XU1288 n1382 n1383 NETTRAN_DUMMY_7784 NETTRAN_DUMMY_7785 INV_X1 
XU1289 n438 n1384 NETTRAN_DUMMY_7786 NETTRAN_DUMMY_7787 INV_X1 
XU1290 n1381 n1385 NETTRAN_DUMMY_7788 NETTRAN_DUMMY_7789 INV_X32 
XU1291 n1391 n1386 NETTRAN_DUMMY_7790 NETTRAN_DUMMY_7791 INV_X1 
XU1292 n1386 n1387 NETTRAN_DUMMY_7792 NETTRAN_DUMMY_7793 INV_X32 
XU1293 n1390 n1388 NETTRAN_DUMMY_7794 NETTRAN_DUMMY_7795 INV_X32 
XU1294 n1388 n1389 NETTRAN_DUMMY_7796 NETTRAN_DUMMY_7797 INV_X1 
XU1295 n433 n1390 NETTRAN_DUMMY_7798 NETTRAN_DUMMY_7799 INV_X1 
XU1296 n1389 n1391 NETTRAN_DUMMY_7800 NETTRAN_DUMMY_7801 INV_X32 
XU1297 n420 n1392 NETTRAN_DUMMY_7802 NETTRAN_DUMMY_7803 INV_X1 
XU1298 n1392 n1393 NETTRAN_DUMMY_7804 NETTRAN_DUMMY_7805 INV_X32 
XU1299 n1393 n1394 NETTRAN_DUMMY_7806 NETTRAN_DUMMY_7807 INV_X1 
XU1300 n1394 n1395 NETTRAN_DUMMY_7808 NETTRAN_DUMMY_7809 INV_X32 
XU1301 n171 n1396 NETTRAN_DUMMY_7810 NETTRAN_DUMMY_7811 CLKBUF_X1 
XU1302 n1398 n1397 NETTRAN_DUMMY_7812 NETTRAN_DUMMY_7813 CLKBUF_X1 
XU1303 n407 n1398 NETTRAN_DUMMY_7814 NETTRAN_DUMMY_7815 INV_X1 
XU1304 n1397 n1399 NETTRAN_DUMMY_7816 NETTRAN_DUMMY_7817 INV_X32 
XU1305 n1399 n1400 NETTRAN_DUMMY_7818 NETTRAN_DUMMY_7819 INV_X1 
XU1306 n1400 n1401 NETTRAN_DUMMY_7820 NETTRAN_DUMMY_7821 INV_X32 
XU1307 n644 n1402 NETTRAN_DUMMY_7822 NETTRAN_DUMMY_7823 INV_X32 
XU1308 n1402 n1403 NETTRAN_DUMMY_7824 NETTRAN_DUMMY_7825 INV_X1 
XU1309 n394 n1404 NETTRAN_DUMMY_7826 NETTRAN_DUMMY_7827 INV_X1 
XU1310 n1403 n1405 NETTRAN_DUMMY_7828 NETTRAN_DUMMY_7829 INV_X32 
XU1311 n145 n1406 NETTRAN_DUMMY_7830 NETTRAN_DUMMY_7831 BUF_X1 
XU1312 n1410 n1407 NETTRAN_DUMMY_7832 NETTRAN_DUMMY_7833 CLKBUF_X1 
XU1313 n1407 n1408 NETTRAN_DUMMY_7834 NETTRAN_DUMMY_7835 INV_X32 
XU1314 n1408 n1409 NETTRAN_DUMMY_7836 NETTRAN_DUMMY_7837 INV_X1 
XU1315 n381 n1410 NETTRAN_DUMMY_7838 NETTRAN_DUMMY_7839 INV_X1 
XU1316 n1409 n1411 NETTRAN_DUMMY_7840 NETTRAN_DUMMY_7841 INV_X32 
XU1317 n1416 n1412 NETTRAN_DUMMY_7842 NETTRAN_DUMMY_7843 BUF_X1 
XU1318 n1415 n1413 NETTRAN_DUMMY_7844 NETTRAN_DUMMY_7845 INV_X32 
XU1319 n1413 n1414 NETTRAN_DUMMY_7846 NETTRAN_DUMMY_7847 INV_X1 
XU1320 n426 n1415 NETTRAN_DUMMY_7848 NETTRAN_DUMMY_7849 INV_X1 
XU1321 n1414 n1416 NETTRAN_DUMMY_7850 NETTRAN_DUMMY_7851 INV_X32 
XU1322 n177 n1417 NETTRAN_DUMMY_7852 NETTRAN_DUMMY_7853 INV_X1 
XU1323 n1417 n1418 NETTRAN_DUMMY_7854 NETTRAN_DUMMY_7855 INV_X32 
XU1324 n413 n1419 NETTRAN_DUMMY_7856 NETTRAN_DUMMY_7857 INV_X1 
XU1325 n1419 n1420 NETTRAN_DUMMY_7858 NETTRAN_DUMMY_7859 INV_X32 
XU1326 n1420 n1421 NETTRAN_DUMMY_7860 NETTRAN_DUMMY_7861 INV_X1 
XU1327 n1421 n1422 NETTRAN_DUMMY_7862 NETTRAN_DUMMY_7863 INV_X32 
XU1328 n1424 n1423 NETTRAN_DUMMY_7864 NETTRAN_DUMMY_7865 CLKBUF_X1 
XU1329 n400 n1424 NETTRAN_DUMMY_7866 NETTRAN_DUMMY_7867 INV_X1 
XU1330 n1423 n1425 NETTRAN_DUMMY_7868 NETTRAN_DUMMY_7869 INV_X32 
XU1331 n1425 n1426 NETTRAN_DUMMY_7870 NETTRAN_DUMMY_7871 INV_X1 
XU1332 n1426 n1427 NETTRAN_DUMMY_7872 NETTRAN_DUMMY_7873 INV_X32 
XU1333 n1429 n1428 NETTRAN_DUMMY_7874 NETTRAN_DUMMY_7875 CLKBUF_X1 
XU1334 n387 n1429 NETTRAN_DUMMY_7876 NETTRAN_DUMMY_7877 INV_X1 
XU1335 n1428 n1430 NETTRAN_DUMMY_7878 NETTRAN_DUMMY_7879 INV_X32 
XU1336 n1430 n1431 NETTRAN_DUMMY_7880 NETTRAN_DUMMY_7881 INV_X1 
XU1337 n1431 n1432 NETTRAN_DUMMY_7882 NETTRAN_DUMMY_7883 INV_X32 
XU1338 n1436 n1433 NETTRAN_DUMMY_7884 NETTRAN_DUMMY_7885 CLKBUF_X1 
XU1339 n1433 n1434 NETTRAN_DUMMY_7886 NETTRAN_DUMMY_7887 INV_X32 
XU1340 n1434 n1435 NETTRAN_DUMMY_7888 NETTRAN_DUMMY_7889 INV_X1 
XU1341 n432 n1436 NETTRAN_DUMMY_7890 NETTRAN_DUMMY_7891 INV_X1 
XU1342 n1435 n1437 NETTRAN_DUMMY_7892 NETTRAN_DUMMY_7893 INV_X32 
XU1343 n1443 n1438 NETTRAN_DUMMY_7894 NETTRAN_DUMMY_7895 INV_X1 
XU1344 n1438 n1439 NETTRAN_DUMMY_7896 NETTRAN_DUMMY_7897 INV_X32 
XU1345 n1442 n1440 NETTRAN_DUMMY_7898 NETTRAN_DUMMY_7899 INV_X32 
XU1346 n1440 n1441 NETTRAN_DUMMY_7900 NETTRAN_DUMMY_7901 INV_X1 
XU1347 n419 n1442 NETTRAN_DUMMY_7902 NETTRAN_DUMMY_7903 INV_X1 
XU1348 n1441 n1443 NETTRAN_DUMMY_7904 NETTRAN_DUMMY_7905 INV_X32 
XU1349 n1447 n1444 NETTRAN_DUMMY_7906 NETTRAN_DUMMY_7907 CLKBUF_X1 
XU1350 n1444 n1445 NETTRAN_DUMMY_7908 NETTRAN_DUMMY_7909 INV_X32 
XU1351 n1445 n1446 NETTRAN_DUMMY_7910 NETTRAN_DUMMY_7911 INV_X1 
XU1352 n406 n1447 NETTRAN_DUMMY_7912 NETTRAN_DUMMY_7913 INV_X1 
XU1353 n1446 n1448 NETTRAN_DUMMY_7914 NETTRAN_DUMMY_7915 INV_X32 
XU1354 n1454 n1449 NETTRAN_DUMMY_7916 NETTRAN_DUMMY_7917 INV_X1 
XU1355 n1449 n1450 NETTRAN_DUMMY_7918 NETTRAN_DUMMY_7919 INV_X32 
XU1356 n393 n1451 NETTRAN_DUMMY_7920 NETTRAN_DUMMY_7921 INV_X1 
XU1357 n1451 n1452 NETTRAN_DUMMY_7922 NETTRAN_DUMMY_7923 INV_X32 
XU1358 n1452 n1453 NETTRAN_DUMMY_7924 NETTRAN_DUMMY_7925 INV_X1 
XU1359 n1453 n1454 NETTRAN_DUMMY_7926 NETTRAN_DUMMY_7927 INV_X32 
XU1360 n1458 n1455 NETTRAN_DUMMY_7928 NETTRAN_DUMMY_7929 CLKBUF_X1 
XU1361 n1455 n1456 NETTRAN_DUMMY_7930 NETTRAN_DUMMY_7931 INV_X32 
XU1362 n1456 n1457 NETTRAN_DUMMY_7932 NETTRAN_DUMMY_7933 INV_X1 
XU1363 n380 n1458 NETTRAN_DUMMY_7934 NETTRAN_DUMMY_7935 INV_X1 
XU1364 n1457 n1459 NETTRAN_DUMMY_7936 NETTRAN_DUMMY_7937 INV_X32 
XU1365 n1465 n1460 NETTRAN_DUMMY_7938 NETTRAN_DUMMY_7939 INV_X1 
XU1366 n1460 n1461 NETTRAN_DUMMY_7940 NETTRAN_DUMMY_7941 INV_X32 
XU1367 n1464 n1462 NETTRAN_DUMMY_7942 NETTRAN_DUMMY_7943 INV_X32 
XU1368 n1462 n1463 NETTRAN_DUMMY_7944 NETTRAN_DUMMY_7945 INV_X1 
XU1369 n425 n1464 NETTRAN_DUMMY_7946 NETTRAN_DUMMY_7947 INV_X1 
XU1370 n1463 n1465 NETTRAN_DUMMY_7948 NETTRAN_DUMMY_7949 INV_X32 
XU1371 n652 n1466 NETTRAN_DUMMY_7950 NETTRAN_DUMMY_7951 INV_X32 
XU1372 n1466 n1467 NETTRAN_DUMMY_7952 NETTRAN_DUMMY_7953 INV_X1 
XU1373 n412 n1468 NETTRAN_DUMMY_7954 NETTRAN_DUMMY_7955 INV_X1 
XU1374 n1467 n1469 NETTRAN_DUMMY_7956 NETTRAN_DUMMY_7957 INV_X32 
XU1375 n163 n1470 NETTRAN_DUMMY_7958 NETTRAN_DUMMY_7959 CLKBUF_X1 
XU1376 n1474 n1471 NETTRAN_DUMMY_7960 NETTRAN_DUMMY_7961 CLKBUF_X1 
XU1377 n1471 n1472 NETTRAN_DUMMY_7962 NETTRAN_DUMMY_7963 INV_X32 
XU1378 n1472 n1473 NETTRAN_DUMMY_7964 NETTRAN_DUMMY_7965 INV_X1 
XU1379 n399 n1474 NETTRAN_DUMMY_7966 NETTRAN_DUMMY_7967 INV_X1 
XU1380 n1473 n1475 NETTRAN_DUMMY_7968 NETTRAN_DUMMY_7969 INV_X32 
XU1381 n1477 n1476 NETTRAN_DUMMY_7970 NETTRAN_DUMMY_7971 CLKBUF_X1 
XU1382 n386 n1477 NETTRAN_DUMMY_7972 NETTRAN_DUMMY_7973 INV_X1 
XU1383 n1476 n1478 NETTRAN_DUMMY_7974 NETTRAN_DUMMY_7975 INV_X32 
XU1384 n1478 n1479 NETTRAN_DUMMY_7976 NETTRAN_DUMMY_7977 INV_X1 
XU1385 n1479 n1480 NETTRAN_DUMMY_7978 NETTRAN_DUMMY_7979 INV_X32 
XU1386 n1486 n1481 NETTRAN_DUMMY_7980 NETTRAN_DUMMY_7981 INV_X1 
XU1387 n1481 n1482 NETTRAN_DUMMY_7982 NETTRAN_DUMMY_7983 INV_X32 
XU1388 n431 n1483 NETTRAN_DUMMY_7984 NETTRAN_DUMMY_7985 INV_X1 
XU1389 n1483 n1484 NETTRAN_DUMMY_7986 NETTRAN_DUMMY_7987 INV_X32 
XU1390 n1484 n1485 NETTRAN_DUMMY_7988 NETTRAN_DUMMY_7989 INV_X1 
XU1391 n1485 n1486 NETTRAN_DUMMY_7990 NETTRAN_DUMMY_7991 INV_X32 
XU1392 n1490 n1487 NETTRAN_DUMMY_7992 NETTRAN_DUMMY_7993 INV_X1 
XU1393 n1487 n1488 NETTRAN_DUMMY_7994 NETTRAN_DUMMY_7995 INV_X32 
XU1394 n418 n1489 NETTRAN_DUMMY_7996 NETTRAN_DUMMY_7997 INV_X1 
XU1395 n1489 n1490 NETTRAN_DUMMY_7998 NETTRAN_DUMMY_7999 INV_X32 
XU1396 n169 n1491 NETTRAN_DUMMY_8000 NETTRAN_DUMMY_8001 BUF_X1 
XU1397 n1493 n1492 NETTRAN_DUMMY_8002 NETTRAN_DUMMY_8003 CLKBUF_X1 
XU1398 n405 n1493 NETTRAN_DUMMY_8004 NETTRAN_DUMMY_8005 INV_X1 
XU1399 n1492 n1494 NETTRAN_DUMMY_8006 NETTRAN_DUMMY_8007 INV_X32 
XU1400 n1494 n1495 NETTRAN_DUMMY_8008 NETTRAN_DUMMY_8009 INV_X1 
XU1401 n1495 n1496 NETTRAN_DUMMY_8010 NETTRAN_DUMMY_8011 INV_X32 
XU1402 n1500 n1497 NETTRAN_DUMMY_8012 NETTRAN_DUMMY_8013 CLKBUF_X1 
XU1403 n392 n1498 NETTRAN_DUMMY_8014 NETTRAN_DUMMY_8015 INV_X1 
XU1404 n1498 n1499 NETTRAN_DUMMY_8016 NETTRAN_DUMMY_8017 INV_X32 
XU1405 n1499 n1500 NETTRAN_DUMMY_8018 NETTRAN_DUMMY_8019 INV_X1 
XU1406 n1497 n1501 NETTRAN_DUMMY_8020 NETTRAN_DUMMY_8021 INV_X32 
XU1407 n1505 n1502 NETTRAN_DUMMY_8022 NETTRAN_DUMMY_8023 CLKBUF_X1 
XU1408 n1502 n1503 NETTRAN_DUMMY_8024 NETTRAN_DUMMY_8025 INV_X32 
XU1409 n1503 n1504 NETTRAN_DUMMY_8026 NETTRAN_DUMMY_8027 INV_X1 
XU1410 n379 n1505 NETTRAN_DUMMY_8028 NETTRAN_DUMMY_8029 INV_X1 
XU1411 n1504 n1506 NETTRAN_DUMMY_8030 NETTRAN_DUMMY_8031 INV_X32 
XU1412 n1510 n1507 NETTRAN_DUMMY_8032 NETTRAN_DUMMY_8033 CLKBUF_X1 
XU1413 n1507 n1508 NETTRAN_DUMMY_8034 NETTRAN_DUMMY_8035 INV_X32 
XU1414 n1508 n1509 NETTRAN_DUMMY_8036 NETTRAN_DUMMY_8037 INV_X1 
XU1415 n424 n1510 NETTRAN_DUMMY_8038 NETTRAN_DUMMY_8039 INV_X1 
XU1416 n1509 n1511 NETTRAN_DUMMY_8040 NETTRAN_DUMMY_8041 INV_X32 
XU1417 n1513 n1512 NETTRAN_DUMMY_8042 NETTRAN_DUMMY_8043 CLKBUF_X1 
XU1418 n411 n1513 NETTRAN_DUMMY_8044 NETTRAN_DUMMY_8045 INV_X1 
XU1419 n1512 n1514 NETTRAN_DUMMY_8046 NETTRAN_DUMMY_8047 INV_X32 
XU1420 n1514 n1515 NETTRAN_DUMMY_8048 NETTRAN_DUMMY_8049 INV_X1 
XU1421 n1515 n1516 NETTRAN_DUMMY_8050 NETTRAN_DUMMY_8051 INV_X32 
XU1422 n1520 n1517 NETTRAN_DUMMY_8052 NETTRAN_DUMMY_8053 CLKBUF_X1 
XU1423 n1517 n1518 NETTRAN_DUMMY_8054 NETTRAN_DUMMY_8055 INV_X32 
XU1424 n1518 n1519 NETTRAN_DUMMY_8056 NETTRAN_DUMMY_8057 INV_X1 
XU1425 n398 n1520 NETTRAN_DUMMY_8058 NETTRAN_DUMMY_8059 INV_X1 
XU1426 n1519 n1521 NETTRAN_DUMMY_8060 NETTRAN_DUMMY_8061 INV_X32 
XU1427 n1525 n1522 NETTRAN_DUMMY_8062 NETTRAN_DUMMY_8063 CLKBUF_X1 
XU1428 n1522 n1523 NETTRAN_DUMMY_8064 NETTRAN_DUMMY_8065 INV_X32 
XU1429 n1523 n1524 NETTRAN_DUMMY_8066 NETTRAN_DUMMY_8067 INV_X1 
XU1430 n385 n1525 NETTRAN_DUMMY_8068 NETTRAN_DUMMY_8069 INV_X1 
XU1431 n1524 n1526 NETTRAN_DUMMY_8070 NETTRAN_DUMMY_8071 INV_X32 
XU1432 n1530 n1527 NETTRAN_DUMMY_8072 NETTRAN_DUMMY_8073 CLKBUF_X1 
XU1433 n1527 n1528 NETTRAN_DUMMY_8074 NETTRAN_DUMMY_8075 INV_X32 
XU1434 n1528 n1529 NETTRAN_DUMMY_8076 NETTRAN_DUMMY_8077 INV_X1 
XU1435 n430 n1530 NETTRAN_DUMMY_8078 NETTRAN_DUMMY_8079 INV_X1 
XU1436 n1529 n1531 NETTRAN_DUMMY_8080 NETTRAN_DUMMY_8081 INV_X32 
XU1437 n417 n1532 NETTRAN_DUMMY_8082 NETTRAN_DUMMY_8083 INV_X1 
XU1438 n1532 n1533 NETTRAN_DUMMY_8084 NETTRAN_DUMMY_8085 INV_X32 
XU1439 n1533 n1534 NETTRAN_DUMMY_8086 NETTRAN_DUMMY_8087 INV_X1 
XU1440 n1534 n1535 NETTRAN_DUMMY_8088 NETTRAN_DUMMY_8089 INV_X32 
XU1441 n168 n1536 NETTRAN_DUMMY_8090 NETTRAN_DUMMY_8091 INV_X1 
XU1442 n1536 n1537 NETTRAN_DUMMY_8092 NETTRAN_DUMMY_8093 INV_X32 
XU1443 n1539 n1538 NETTRAN_DUMMY_8094 NETTRAN_DUMMY_8095 CLKBUF_X1 
XU1444 n404 n1539 NETTRAN_DUMMY_8096 NETTRAN_DUMMY_8097 INV_X1 
XU1445 n1538 n1540 NETTRAN_DUMMY_8098 NETTRAN_DUMMY_8099 INV_X32 
XU1446 n1540 n1541 NETTRAN_DUMMY_8100 NETTRAN_DUMMY_8101 INV_X1 
XU1447 n1541 n1542 NETTRAN_DUMMY_8102 NETTRAN_DUMMY_8103 INV_X32 
XU1448 n1546 n1543 NETTRAN_DUMMY_8104 NETTRAN_DUMMY_8105 CLKBUF_X1 
XU1449 n391 n1544 NETTRAN_DUMMY_8106 NETTRAN_DUMMY_8107 INV_X1 
XU1450 n1544 n1545 NETTRAN_DUMMY_8108 NETTRAN_DUMMY_8109 INV_X32 
XU1451 n1545 n1546 NETTRAN_DUMMY_8110 NETTRAN_DUMMY_8111 INV_X1 
XU1452 n1543 n1547 NETTRAN_DUMMY_8112 NETTRAN_DUMMY_8113 INV_X32 
XU1453 n1551 n1548 NETTRAN_DUMMY_8114 NETTRAN_DUMMY_8115 CLKBUF_X1 
XU1454 n1548 n1549 NETTRAN_DUMMY_8116 NETTRAN_DUMMY_8117 INV_X32 
XU1455 n1549 n1550 NETTRAN_DUMMY_8118 NETTRAN_DUMMY_8119 INV_X1 
XU1456 n378 n1551 NETTRAN_DUMMY_8120 NETTRAN_DUMMY_8121 INV_X1 
XU1457 n1550 n1552 NETTRAN_DUMMY_8122 NETTRAN_DUMMY_8123 INV_X32 
XU1458 n1558 n1553 NETTRAN_DUMMY_8124 NETTRAN_DUMMY_8125 INV_X1 
XU1459 n1553 n1554 NETTRAN_DUMMY_8126 NETTRAN_DUMMY_8127 INV_X32 
XU1460 n1557 n1555 NETTRAN_DUMMY_8128 NETTRAN_DUMMY_8129 INV_X32 
XU1461 n1555 n1556 NETTRAN_DUMMY_8130 NETTRAN_DUMMY_8131 INV_X1 
XU1462 n423 n1557 NETTRAN_DUMMY_8132 NETTRAN_DUMMY_8133 INV_X1 
XU1463 n1556 n1558 NETTRAN_DUMMY_8134 NETTRAN_DUMMY_8135 INV_X32 
XU1464 n1564 n1559 NETTRAN_DUMMY_8136 NETTRAN_DUMMY_8137 INV_X1 
XU1465 n1559 n1560 NETTRAN_DUMMY_8138 NETTRAN_DUMMY_8139 INV_X32 
XU1466 n410 n1561 NETTRAN_DUMMY_8140 NETTRAN_DUMMY_8141 INV_X1 
XU1467 n1561 n1562 NETTRAN_DUMMY_8142 NETTRAN_DUMMY_8143 INV_X32 
XU1468 n1562 n1563 NETTRAN_DUMMY_8144 NETTRAN_DUMMY_8145 INV_X1 
XU1469 n1563 n1564 NETTRAN_DUMMY_8146 NETTRAN_DUMMY_8147 INV_X32 
XU1470 n1569 n1565 NETTRAN_DUMMY_8148 NETTRAN_DUMMY_8149 BUF_X1 
XU1471 n1568 n1566 NETTRAN_DUMMY_8150 NETTRAN_DUMMY_8151 INV_X32 
XU1472 n1566 n1567 NETTRAN_DUMMY_8152 NETTRAN_DUMMY_8153 INV_X1 
XU1473 n397 n1568 NETTRAN_DUMMY_8154 NETTRAN_DUMMY_8155 INV_X1 
XU1474 n1567 n1569 NETTRAN_DUMMY_8156 NETTRAN_DUMMY_8157 INV_X32 
XU1475 n673 n1570 NETTRAN_DUMMY_8158 NETTRAN_DUMMY_8159 INV_X32 
XU1476 n1570 n1571 NETTRAN_DUMMY_8160 NETTRAN_DUMMY_8161 INV_X1 
XU1477 n1572 n1573 NETTRAN_DUMMY_8162 NETTRAN_DUMMY_8163 INV_X1 
XU1478 n384 n1574 NETTRAN_DUMMY_8164 NETTRAN_DUMMY_8165 INV_X1 
XU1479 n1571 n1575 NETTRAN_DUMMY_8166 NETTRAN_DUMMY_8167 INV_X32 
XU1480 n1579 n1576 NETTRAN_DUMMY_8168 NETTRAN_DUMMY_8169 INV_X1 
XU1481 n1576 n1577 NETTRAN_DUMMY_8170 NETTRAN_DUMMY_8171 INV_X32 
XU1482 n429 n1578 NETTRAN_DUMMY_8172 NETTRAN_DUMMY_8173 INV_X1 
XU1483 n1578 n1579 NETTRAN_DUMMY_8174 NETTRAN_DUMMY_8175 INV_X32 
XU1484 n180 n1580 NETTRAN_DUMMY_8176 NETTRAN_DUMMY_8177 INV_X32 
XU1485 n1580 n1581 NETTRAN_DUMMY_8178 NETTRAN_DUMMY_8179 INV_X1 
XU1486 n1586 n1582 NETTRAN_DUMMY_8180 NETTRAN_DUMMY_8181 INV_X32 
XU1487 n1582 n1583 NETTRAN_DUMMY_8182 NETTRAN_DUMMY_8183 INV_X1 
XU1488 n1583 n1584 NETTRAN_DUMMY_8184 NETTRAN_DUMMY_8185 INV_X32 
XU1489 n1584 n1585 NETTRAN_DUMMY_8186 NETTRAN_DUMMY_8187 INV_X1 
XU1490 n416 n1586 NETTRAN_DUMMY_8188 NETTRAN_DUMMY_8189 INV_X1 
XU1491 n1585 n1587 NETTRAN_DUMMY_8190 NETTRAN_DUMMY_8191 INV_X32 
XU1492 n1589 n1588 NETTRAN_DUMMY_8192 NETTRAN_DUMMY_8193 CLKBUF_X1 
XU1493 n403 n1589 NETTRAN_DUMMY_8194 NETTRAN_DUMMY_8195 INV_X1 
XU1494 n1588 n1590 NETTRAN_DUMMY_8196 NETTRAN_DUMMY_8197 INV_X32 
XU1495 n1590 n1591 NETTRAN_DUMMY_8198 NETTRAN_DUMMY_8199 INV_X1 
XU1496 n1591 n1592 NETTRAN_DUMMY_8200 NETTRAN_DUMMY_8201 INV_X32 
XU1497 n1596 n1593 NETTRAN_DUMMY_8202 NETTRAN_DUMMY_8203 CLKBUF_X1 
XU1498 n1593 n1594 NETTRAN_DUMMY_8204 NETTRAN_DUMMY_8205 INV_X32 
XU1499 n1594 n1595 NETTRAN_DUMMY_8206 NETTRAN_DUMMY_8207 INV_X1 
XU1500 n390 n1596 NETTRAN_DUMMY_8208 NETTRAN_DUMMY_8209 INV_X1 
XU1501 n1595 n1597 NETTRAN_DUMMY_8210 NETTRAN_DUMMY_8211 INV_X32 
XU1502 n1601 n1598 NETTRAN_DUMMY_8212 NETTRAN_DUMMY_8213 CLKBUF_X1 
XU1503 n1598 n1599 NETTRAN_DUMMY_8214 NETTRAN_DUMMY_8215 INV_X32 
XU1504 n1599 n1600 NETTRAN_DUMMY_8216 NETTRAN_DUMMY_8217 INV_X1 
XU1505 n377 n1601 NETTRAN_DUMMY_8218 NETTRAN_DUMMY_8219 INV_X1 
XU1506 n1600 n1602 NETTRAN_DUMMY_8220 NETTRAN_DUMMY_8221 INV_X32 
XU1507 n1608 n1603 NETTRAN_DUMMY_8222 NETTRAN_DUMMY_8223 INV_X1 
XU1508 n1603 n1604 NETTRAN_DUMMY_8224 NETTRAN_DUMMY_8225 INV_X32 
XU1509 n1607 n1605 NETTRAN_DUMMY_8226 NETTRAN_DUMMY_8227 INV_X32 
XU1510 n1605 n1606 NETTRAN_DUMMY_8228 NETTRAN_DUMMY_8229 INV_X1 
XU1511 n422 n1607 NETTRAN_DUMMY_8230 NETTRAN_DUMMY_8231 INV_X1 
XU1512 n1606 n1608 NETTRAN_DUMMY_8232 NETTRAN_DUMMY_8233 INV_X32 
XU1513 n1610 n1609 NETTRAN_DUMMY_8234 NETTRAN_DUMMY_8235 CLKBUF_X1 
XU1514 n1613 n1610 NETTRAN_DUMMY_8236 NETTRAN_DUMMY_8237 INV_X1 
XU1515 n1609 n1611 NETTRAN_DUMMY_8238 NETTRAN_DUMMY_8239 INV_X32 
XU1516 n409 n1612 NETTRAN_DUMMY_8240 NETTRAN_DUMMY_8241 INV_X1 
XU1517 n1612 n1613 NETTRAN_DUMMY_8242 NETTRAN_DUMMY_8243 INV_X32 
XU1518 n1617 n1614 NETTRAN_DUMMY_8244 NETTRAN_DUMMY_8245 CLKBUF_X1 
XU1519 n1614 n1615 NETTRAN_DUMMY_8246 NETTRAN_DUMMY_8247 INV_X32 
XU1520 n1615 n1616 NETTRAN_DUMMY_8248 NETTRAN_DUMMY_8249 INV_X1 
XU1521 n396 n1617 NETTRAN_DUMMY_8250 NETTRAN_DUMMY_8251 INV_X1 
XU1522 n1616 n1618 NETTRAN_DUMMY_8252 NETTRAN_DUMMY_8253 INV_X32 
XU1523 n1622 n1619 NETTRAN_DUMMY_8254 NETTRAN_DUMMY_8255 CLKBUF_X1 
XU1524 n383 n1620 NETTRAN_DUMMY_8256 NETTRAN_DUMMY_8257 INV_X1 
XU1525 n1620 n1621 NETTRAN_DUMMY_8258 NETTRAN_DUMMY_8259 INV_X32 
XU1526 n1621 n1622 NETTRAN_DUMMY_8260 NETTRAN_DUMMY_8261 INV_X1 
XU1527 n1619 n1623 NETTRAN_DUMMY_8262 NETTRAN_DUMMY_8263 INV_X32 
XU1528 n1629 n1624 NETTRAN_DUMMY_8264 NETTRAN_DUMMY_8265 INV_X1 
XU1529 n1624 n1625 NETTRAN_DUMMY_8266 NETTRAN_DUMMY_8267 INV_X32 
XU1530 n1628 n1626 NETTRAN_DUMMY_8268 NETTRAN_DUMMY_8269 INV_X32 
XU1531 n1626 n1627 NETTRAN_DUMMY_8270 NETTRAN_DUMMY_8271 INV_X1 
XU1532 n428 n1628 NETTRAN_DUMMY_8272 NETTRAN_DUMMY_8273 INV_X1 
XU1533 n1627 n1629 NETTRAN_DUMMY_8274 NETTRAN_DUMMY_8275 INV_X32 
XU1534 n1635 n1630 NETTRAN_DUMMY_8276 NETTRAN_DUMMY_8277 INV_X1 
XU1535 n1630 n1631 NETTRAN_DUMMY_8278 NETTRAN_DUMMY_8279 INV_X32 
XU1536 n1634 n1632 NETTRAN_DUMMY_8280 NETTRAN_DUMMY_8281 INV_X32 
XU1537 n1632 n1633 NETTRAN_DUMMY_8282 NETTRAN_DUMMY_8283 INV_X1 
XU1538 n415 n1634 NETTRAN_DUMMY_8284 NETTRAN_DUMMY_8285 INV_X1 
XU1539 n1633 n1635 NETTRAN_DUMMY_8286 NETTRAN_DUMMY_8287 INV_X32 
XU1540 n682 n1636 NETTRAN_DUMMY_8288 NETTRAN_DUMMY_8289 INV_X32 
XU1541 n1636 n1637 NETTRAN_DUMMY_8290 NETTRAN_DUMMY_8291 INV_X1 
XU1542 n551 n1638 NETTRAN_DUMMY_8292 NETTRAN_DUMMY_8293 INV_X1 
XU1543 n1637 n1639 NETTRAN_DUMMY_8294 NETTRAN_DUMMY_8295 INV_X32 
XU1544 n55 n1640 NETTRAN_DUMMY_8296 NETTRAN_DUMMY_8297 CLKBUF_X1 
XU1545 n1643 n1641 NETTRAN_DUMMY_8298 NETTRAN_DUMMY_8299 INV_X32 
XU1546 n1641 n1642 NETTRAN_DUMMY_8300 NETTRAN_DUMMY_8301 INV_X1 
XU1547 n544 n1643 NETTRAN_DUMMY_8302 NETTRAN_DUMMY_8303 INV_X1 
XU1548 n1642 n1644 NETTRAN_DUMMY_8304 NETTRAN_DUMMY_8305 INV_X32 
XU1549 n48 n1645 NETTRAN_DUMMY_8306 NETTRAN_DUMMY_8307 INV_X1 
XU1550 n1645 n1646 NETTRAN_DUMMY_8308 NETTRAN_DUMMY_8309 INV_X32 
XU1551 n1648 n1647 NETTRAN_DUMMY_8310 NETTRAN_DUMMY_8311 CLKBUF_X1 
XU1552 n537 n1648 NETTRAN_DUMMY_8312 NETTRAN_DUMMY_8313 INV_X1 
XU1553 n1647 n1649 NETTRAN_DUMMY_8314 NETTRAN_DUMMY_8315 INV_X32 
XU1554 n1649 n1650 NETTRAN_DUMMY_8316 NETTRAN_DUMMY_8317 INV_X1 
XU1555 n1650 n1651 NETTRAN_DUMMY_8318 NETTRAN_DUMMY_8319 INV_X32 
XU1556 n1655 n1652 NETTRAN_DUMMY_8320 NETTRAN_DUMMY_8321 CLKBUF_X1 
XU1557 n1652 n1653 NETTRAN_DUMMY_8322 NETTRAN_DUMMY_8323 INV_X32 
XU1558 n1653 n1654 NETTRAN_DUMMY_8324 NETTRAN_DUMMY_8325 INV_X1 
XU1559 n530 n1655 NETTRAN_DUMMY_8326 NETTRAN_DUMMY_8327 INV_X1 
XU1560 n1654 n1656 NETTRAN_DUMMY_8328 NETTRAN_DUMMY_8329 INV_X32 
XU1561 n1658 n1657 NETTRAN_DUMMY_8330 NETTRAN_DUMMY_8331 CLKBUF_X1 
XU1562 n523 n1658 NETTRAN_DUMMY_8332 NETTRAN_DUMMY_8333 INV_X1 
XU1563 n1657 n1659 NETTRAN_DUMMY_8334 NETTRAN_DUMMY_8335 INV_X32 
XU1564 n1659 n1660 NETTRAN_DUMMY_8336 NETTRAN_DUMMY_8337 INV_X1 
XU1565 n1660 n1661 NETTRAN_DUMMY_8338 NETTRAN_DUMMY_8339 INV_X32 
XU1566 n1663 n1662 NETTRAN_DUMMY_8340 NETTRAN_DUMMY_8341 CLKBUF_X1 
XU1567 n516 n1663 NETTRAN_DUMMY_8342 NETTRAN_DUMMY_8343 INV_X1 
XU1568 n1662 n1664 NETTRAN_DUMMY_8344 NETTRAN_DUMMY_8345 INV_X32 
XU1569 n1664 n1665 NETTRAN_DUMMY_8346 NETTRAN_DUMMY_8347 INV_X1 
XU1570 n1665 n1666 NETTRAN_DUMMY_8348 NETTRAN_DUMMY_8349 INV_X32 
XU1571 n1670 n1667 NETTRAN_DUMMY_8350 NETTRAN_DUMMY_8351 CLKBUF_X1 
XU1572 n1667 n1668 NETTRAN_DUMMY_8352 NETTRAN_DUMMY_8353 INV_X32 
XU1573 n1668 n1669 NETTRAN_DUMMY_8354 NETTRAN_DUMMY_8355 INV_X1 
XU1574 n509 n1670 NETTRAN_DUMMY_8356 NETTRAN_DUMMY_8357 INV_X1 
XU1575 n1669 n1671 NETTRAN_DUMMY_8358 NETTRAN_DUMMY_8359 INV_X32 
XU1576 n689 n1672 NETTRAN_DUMMY_8360 NETTRAN_DUMMY_8361 INV_X32 
XU1577 n1672 n1673 NETTRAN_DUMMY_8362 NETTRAN_DUMMY_8363 INV_X1 
XU1578 n502 n1674 NETTRAN_DUMMY_8364 NETTRAN_DUMMY_8365 INV_X1 
XU1579 n1673 n1675 NETTRAN_DUMMY_8366 NETTRAN_DUMMY_8367 INV_X32 
XU1580 n6 n1676 NETTRAN_DUMMY_8368 NETTRAN_DUMMY_8369 BUF_X1 
XU1581 n1680 n1677 NETTRAN_DUMMY_8370 NETTRAN_DUMMY_8371 INV_X1 
XU1582 n691 n1678 NETTRAN_DUMMY_8372 NETTRAN_DUMMY_8373 INV_X32 
XU1583 n547 n1679 NETTRAN_DUMMY_8374 NETTRAN_DUMMY_8375 INV_X1 
XU1584 n1679 n1680 NETTRAN_DUMMY_8376 NETTRAN_DUMMY_8377 INV_X32 
XU1585 n51 n1681 NETTRAN_DUMMY_8378 NETTRAN_DUMMY_8379 BUF_X1 
XU1586 n1683 n1682 NETTRAN_DUMMY_8380 NETTRAN_DUMMY_8381 CLKBUF_X1 
XU1587 n540 n1683 NETTRAN_DUMMY_8382 NETTRAN_DUMMY_8383 INV_X1 
XU1588 n1682 n1684 NETTRAN_DUMMY_8384 NETTRAN_DUMMY_8385 INV_X32 
XU1589 n1684 n1685 NETTRAN_DUMMY_8386 NETTRAN_DUMMY_8387 INV_X1 
XU1590 n1685 n1686 NETTRAN_DUMMY_8388 NETTRAN_DUMMY_8389 INV_X32 
XU1591 n1692 n1687 NETTRAN_DUMMY_8390 NETTRAN_DUMMY_8391 INV_X1 
XU1592 n1687 n1688 NETTRAN_DUMMY_8392 NETTRAN_DUMMY_8393 INV_X32 
XU1593 n1691 n1689 NETTRAN_DUMMY_8394 NETTRAN_DUMMY_8395 INV_X32 
XU1594 n1689 n1690 NETTRAN_DUMMY_8396 NETTRAN_DUMMY_8397 INV_X1 
XU1595 n533 n1691 NETTRAN_DUMMY_8398 NETTRAN_DUMMY_8399 INV_X1 
XU1596 n1690 n1692 NETTRAN_DUMMY_8400 NETTRAN_DUMMY_8401 INV_X32 
XU1597 n1694 n1693 NETTRAN_DUMMY_8402 NETTRAN_DUMMY_8403 CLKBUF_X1 
XU1598 n526 n1694 NETTRAN_DUMMY_8404 NETTRAN_DUMMY_8405 INV_X1 
XU1599 n1693 n1695 NETTRAN_DUMMY_8406 NETTRAN_DUMMY_8407 INV_X32 
XU1600 n1695 n1696 NETTRAN_DUMMY_8408 NETTRAN_DUMMY_8409 INV_X1 
XU1601 n1696 n1697 NETTRAN_DUMMY_8410 NETTRAN_DUMMY_8411 INV_X32 
XU1602 n1701 n1698 NETTRAN_DUMMY_8412 NETTRAN_DUMMY_8413 CLKBUF_X1 
XU1603 n519 n1699 NETTRAN_DUMMY_8414 NETTRAN_DUMMY_8415 INV_X1 
XU1604 n1699 n1700 NETTRAN_DUMMY_8416 NETTRAN_DUMMY_8417 INV_X32 
XU1605 n1700 n1701 NETTRAN_DUMMY_8418 NETTRAN_DUMMY_8419 INV_X1 
XU1606 n1698 n1702 NETTRAN_DUMMY_8420 NETTRAN_DUMMY_8421 INV_X32 
XU1607 n1708 n1703 NETTRAN_DUMMY_8422 NETTRAN_DUMMY_8423 INV_X1 
XU1608 n1703 n1704 NETTRAN_DUMMY_8424 NETTRAN_DUMMY_8425 INV_X32 
XU1609 n512 n1705 NETTRAN_DUMMY_8426 NETTRAN_DUMMY_8427 INV_X1 
XU1610 n1705 n1706 NETTRAN_DUMMY_8428 NETTRAN_DUMMY_8429 INV_X32 
XU1611 n1706 n1707 NETTRAN_DUMMY_8430 NETTRAN_DUMMY_8431 INV_X1 
XU1612 n1707 n1708 NETTRAN_DUMMY_8432 NETTRAN_DUMMY_8433 INV_X32 
XU1613 n1712 n1709 NETTRAN_DUMMY_8434 NETTRAN_DUMMY_8435 CLKBUF_X1 
XU1614 n505 n1710 NETTRAN_DUMMY_8436 NETTRAN_DUMMY_8437 INV_X1 
XU1615 n1710 n1711 NETTRAN_DUMMY_8438 NETTRAN_DUMMY_8439 INV_X32 
XU1616 n1711 n1712 NETTRAN_DUMMY_8440 NETTRAN_DUMMY_8441 INV_X1 
XU1617 n1709 n1713 NETTRAN_DUMMY_8442 NETTRAN_DUMMY_8443 INV_X32 
XU1618 n498 n1714 NETTRAN_DUMMY_8444 NETTRAN_DUMMY_8445 INV_X1 
XU1619 n1714 n1715 NETTRAN_DUMMY_8446 NETTRAN_DUMMY_8447 INV_X32 
XU1620 n1715 n1716 NETTRAN_DUMMY_8448 NETTRAN_DUMMY_8449 INV_X1 
XU1621 n696 n1717 NETTRAN_DUMMY_8450 NETTRAN_DUMMY_8451 INV_X32 
XU1622 n2 n1718 NETTRAN_DUMMY_8452 NETTRAN_DUMMY_8453 INV_X1 
XU1623 n1718 n1719 NETTRAN_DUMMY_8454 NETTRAN_DUMMY_8455 INV_X8 
XU1624 n1723 n1720 NETTRAN_DUMMY_8456 NETTRAN_DUMMY_8457 CLKBUF_X1 
XU1625 n1720 n1721 NETTRAN_DUMMY_8458 NETTRAN_DUMMY_8459 INV_X32 
XU1626 n1721 n1722 NETTRAN_DUMMY_8460 NETTRAN_DUMMY_8461 INV_X1 
XU1627 n550 n1723 NETTRAN_DUMMY_8462 NETTRAN_DUMMY_8463 INV_X1 
XU1628 n1722 n1724 NETTRAN_DUMMY_8464 NETTRAN_DUMMY_8465 INV_X32 
XU1629 n699 n1725 NETTRAN_DUMMY_8466 NETTRAN_DUMMY_8467 INV_X32 
XU1630 n1725 n1726 NETTRAN_DUMMY_8468 NETTRAN_DUMMY_8469 INV_X1 
XU1631 n543 n1727 NETTRAN_DUMMY_8470 NETTRAN_DUMMY_8471 INV_X1 
XU1632 n1726 n1728 NETTRAN_DUMMY_8472 NETTRAN_DUMMY_8473 INV_X32 
XU1633 n47 n1729 NETTRAN_DUMMY_8474 NETTRAN_DUMMY_8475 BUF_X1 
XU1634 n1735 n1730 NETTRAN_DUMMY_8476 NETTRAN_DUMMY_8477 INV_X1 
XU1635 n1730 n1731 NETTRAN_DUMMY_8478 NETTRAN_DUMMY_8479 INV_X32 
XU1636 n1734 n1732 NETTRAN_DUMMY_8480 NETTRAN_DUMMY_8481 INV_X32 
XU1637 n1732 n1733 NETTRAN_DUMMY_8482 NETTRAN_DUMMY_8483 INV_X1 
XU1638 n536 n1734 NETTRAN_DUMMY_8484 NETTRAN_DUMMY_8485 INV_X1 
XU1639 n1733 n1735 NETTRAN_DUMMY_8486 NETTRAN_DUMMY_8487 INV_X32 
XU1640 n1739 n1736 NETTRAN_DUMMY_8488 NETTRAN_DUMMY_8489 CLKBUF_X1 
XU1641 n1736 n1737 NETTRAN_DUMMY_8490 NETTRAN_DUMMY_8491 INV_X32 
XU1642 n1737 n1738 NETTRAN_DUMMY_8492 NETTRAN_DUMMY_8493 INV_X1 
XU1643 n529 n1739 NETTRAN_DUMMY_8494 NETTRAN_DUMMY_8495 INV_X1 
XU1644 n1738 n1740 NETTRAN_DUMMY_8496 NETTRAN_DUMMY_8497 INV_X32 
XU1645 n1744 n1741 NETTRAN_DUMMY_8498 NETTRAN_DUMMY_8499 CLKBUF_X1 
XU1646 n1741 n1742 NETTRAN_DUMMY_8500 NETTRAN_DUMMY_8501 INV_X32 
XU1647 n1742 n1743 NETTRAN_DUMMY_8502 NETTRAN_DUMMY_8503 INV_X1 
XU1648 n522 n1744 NETTRAN_DUMMY_8504 NETTRAN_DUMMY_8505 INV_X1 
XU1649 n1743 n1745 NETTRAN_DUMMY_8506 NETTRAN_DUMMY_8507 INV_X32 
XU1650 n1749 n1746 NETTRAN_DUMMY_8508 NETTRAN_DUMMY_8509 CLKBUF_X1 
XU1651 n1746 n1747 NETTRAN_DUMMY_8510 NETTRAN_DUMMY_8511 INV_X32 
XU1652 n1747 n1748 NETTRAN_DUMMY_8512 NETTRAN_DUMMY_8513 INV_X1 
XU1653 n515 n1749 NETTRAN_DUMMY_8514 NETTRAN_DUMMY_8515 INV_X1 
XU1654 n1748 n1750 NETTRAN_DUMMY_8516 NETTRAN_DUMMY_8517 INV_X32 
XU1655 n1754 n1751 NETTRAN_DUMMY_8518 NETTRAN_DUMMY_8519 CLKBUF_X1 
XU1656 n508 n1752 NETTRAN_DUMMY_8520 NETTRAN_DUMMY_8521 INV_X1 
XU1657 n1752 n1753 NETTRAN_DUMMY_8522 NETTRAN_DUMMY_8523 INV_X32 
XU1658 n1753 n1754 NETTRAN_DUMMY_8524 NETTRAN_DUMMY_8525 INV_X1 
XU1659 n1751 n1755 NETTRAN_DUMMY_8526 NETTRAN_DUMMY_8527 INV_X32 
XU1660 n1757 n1756 NETTRAN_DUMMY_8528 NETTRAN_DUMMY_8529 CLKBUF_X1 
XU1661 n501 n1757 NETTRAN_DUMMY_8530 NETTRAN_DUMMY_8531 INV_X1 
XU1662 n1756 n1758 NETTRAN_DUMMY_8532 NETTRAN_DUMMY_8533 INV_X32 
XU1663 n1758 n1759 NETTRAN_DUMMY_8534 NETTRAN_DUMMY_8535 INV_X1 
XU1664 n1759 n1760 NETTRAN_DUMMY_8536 NETTRAN_DUMMY_8537 INV_X32 
XU1665 n1764 n1761 NETTRAN_DUMMY_8538 NETTRAN_DUMMY_8539 INV_X1 
XU1666 n706 n1762 NETTRAN_DUMMY_8540 NETTRAN_DUMMY_8541 INV_X32 
XU1667 n546 n1763 NETTRAN_DUMMY_8542 NETTRAN_DUMMY_8543 INV_X1 
XU1668 n1763 n1764 NETTRAN_DUMMY_8544 NETTRAN_DUMMY_8545 INV_X32 
XU1669 n50 n1765 NETTRAN_DUMMY_8546 NETTRAN_DUMMY_8547 BUF_X1 
XU1670 n1767 n1766 NETTRAN_DUMMY_8548 NETTRAN_DUMMY_8549 CLKBUF_X1 
XU1671 n539 n1767 NETTRAN_DUMMY_8550 NETTRAN_DUMMY_8551 INV_X1 
XU1672 n1766 n1768 NETTRAN_DUMMY_8552 NETTRAN_DUMMY_8553 INV_X32 
XU1673 n1768 n1769 NETTRAN_DUMMY_8554 NETTRAN_DUMMY_8555 INV_X1 
XU1674 n1769 n1770 NETTRAN_DUMMY_8556 NETTRAN_DUMMY_8557 INV_X32 
XU1675 n1776 n1771 NETTRAN_DUMMY_8558 NETTRAN_DUMMY_8559 INV_X1 
XU1676 n1771 n1772 NETTRAN_DUMMY_8560 NETTRAN_DUMMY_8561 INV_X32 
XU1677 n1775 n1773 NETTRAN_DUMMY_8562 NETTRAN_DUMMY_8563 INV_X32 
XU1678 n1773 n1774 NETTRAN_DUMMY_8564 NETTRAN_DUMMY_8565 INV_X1 
XU1679 n532 n1775 NETTRAN_DUMMY_8566 NETTRAN_DUMMY_8567 INV_X1 
XU1680 n1774 n1776 NETTRAN_DUMMY_8568 NETTRAN_DUMMY_8569 INV_X32 
XU1681 n1780 n1777 NETTRAN_DUMMY_8570 NETTRAN_DUMMY_8571 CLKBUF_X1 
XU1682 n1777 n1778 NETTRAN_DUMMY_8572 NETTRAN_DUMMY_8573 INV_X32 
XU1683 n1778 n1779 NETTRAN_DUMMY_8574 NETTRAN_DUMMY_8575 INV_X1 
XU1684 n525 n1780 NETTRAN_DUMMY_8576 NETTRAN_DUMMY_8577 INV_X1 
XU1685 n1779 n1781 NETTRAN_DUMMY_8578 NETTRAN_DUMMY_8579 INV_X32 
XU1686 n1785 n1782 NETTRAN_DUMMY_8580 NETTRAN_DUMMY_8581 CLKBUF_X1 
XU1687 n518 n1783 NETTRAN_DUMMY_8582 NETTRAN_DUMMY_8583 INV_X1 
XU1688 n1783 n1784 NETTRAN_DUMMY_8584 NETTRAN_DUMMY_8585 INV_X32 
XU1689 n1784 n1785 NETTRAN_DUMMY_8586 NETTRAN_DUMMY_8587 INV_X1 
XU1690 n1782 n1786 NETTRAN_DUMMY_8588 NETTRAN_DUMMY_8589 INV_X32 
XU1691 n1791 n1787 NETTRAN_DUMMY_8590 NETTRAN_DUMMY_8591 BUF_X1 
XU1692 n1790 n1788 NETTRAN_DUMMY_8592 NETTRAN_DUMMY_8593 INV_X32 
XU1693 n1788 n1789 NETTRAN_DUMMY_8594 NETTRAN_DUMMY_8595 INV_X1 
XU1694 n511 n1790 NETTRAN_DUMMY_8596 NETTRAN_DUMMY_8597 INV_X1 
XU1695 n1789 n1791 NETTRAN_DUMMY_8598 NETTRAN_DUMMY_8599 INV_X32 
XU1696 n504 n1792 NETTRAN_DUMMY_8600 NETTRAN_DUMMY_8601 INV_X1 
XU1697 n1792 n1793 NETTRAN_DUMMY_8602 NETTRAN_DUMMY_8603 INV_X32 
XU1698 n1793 n1794 NETTRAN_DUMMY_8604 NETTRAN_DUMMY_8605 INV_X1 
XU1699 n1794 n1795 NETTRAN_DUMMY_8606 NETTRAN_DUMMY_8607 INV_X32 
XU1700 n15 n1796 NETTRAN_DUMMY_8608 NETTRAN_DUMMY_8609 INV_X32 
XU1701 n1796 n1797 NETTRAN_DUMMY_8610 NETTRAN_DUMMY_8611 INV_X1 
XU1702 n1801 n1798 NETTRAN_DUMMY_8612 NETTRAN_DUMMY_8613 CLKBUF_X1 
XU1703 n1798 n1799 NETTRAN_DUMMY_8614 NETTRAN_DUMMY_8615 INV_X32 
XU1704 n1799 n1800 NETTRAN_DUMMY_8616 NETTRAN_DUMMY_8617 INV_X1 
XU1705 n497 n1801 NETTRAN_DUMMY_8618 NETTRAN_DUMMY_8619 INV_X1 
XU1706 n1800 n1802 NETTRAN_DUMMY_8620 NETTRAN_DUMMY_8621 INV_X32 
XU1707 n1808 n1803 NETTRAN_DUMMY_8622 NETTRAN_DUMMY_8623 INV_X1 
XU1708 n1803 n1804 NETTRAN_DUMMY_8624 NETTRAN_DUMMY_8625 INV_X32 
XU1709 n1807 n1805 NETTRAN_DUMMY_8626 NETTRAN_DUMMY_8627 INV_X32 
XU1710 n1805 n1806 NETTRAN_DUMMY_8628 NETTRAN_DUMMY_8629 INV_X1 
XU1711 n549 n1807 NETTRAN_DUMMY_8630 NETTRAN_DUMMY_8631 INV_X1 
XU1712 n1806 n1808 NETTRAN_DUMMY_8632 NETTRAN_DUMMY_8633 INV_X32 
XU1713 n1810 n1809 NETTRAN_DUMMY_8634 NETTRAN_DUMMY_8635 CLKBUF_X1 
XU1714 n542 n1810 NETTRAN_DUMMY_8636 NETTRAN_DUMMY_8637 INV_X1 
XU1715 n1809 n1811 NETTRAN_DUMMY_8638 NETTRAN_DUMMY_8639 INV_X32 
XU1716 n1811 n1812 NETTRAN_DUMMY_8640 NETTRAN_DUMMY_8641 INV_X1 
XU1717 n1812 n1813 NETTRAN_DUMMY_8642 NETTRAN_DUMMY_8643 INV_X32 
XU1718 n1817 n1814 NETTRAN_DUMMY_8644 NETTRAN_DUMMY_8645 CLKBUF_X1 
XU1719 n1814 n1815 NETTRAN_DUMMY_8646 NETTRAN_DUMMY_8647 INV_X32 
XU1720 n1815 n1816 NETTRAN_DUMMY_8648 NETTRAN_DUMMY_8649 INV_X1 
XU1721 n535 n1817 NETTRAN_DUMMY_8650 NETTRAN_DUMMY_8651 INV_X1 
XU1722 n1816 n1818 NETTRAN_DUMMY_8652 NETTRAN_DUMMY_8653 INV_X32 
XU1723 n1822 n1819 NETTRAN_DUMMY_8654 NETTRAN_DUMMY_8655 CLKBUF_X1 
XU1724 n528 n1820 NETTRAN_DUMMY_8656 NETTRAN_DUMMY_8657 INV_X1 
XU1725 n1820 n1821 NETTRAN_DUMMY_8658 NETTRAN_DUMMY_8659 INV_X32 
XU1726 n1821 n1822 NETTRAN_DUMMY_8660 NETTRAN_DUMMY_8661 INV_X1 
XU1727 n1819 n1823 NETTRAN_DUMMY_8662 NETTRAN_DUMMY_8663 INV_X32 
XU1728 n1827 n1824 NETTRAN_DUMMY_8664 NETTRAN_DUMMY_8665 CLKBUF_X1 
XU1729 n1824 n1825 NETTRAN_DUMMY_8666 NETTRAN_DUMMY_8667 INV_X32 
XU1730 n1825 n1826 NETTRAN_DUMMY_8668 NETTRAN_DUMMY_8669 INV_X1 
XU1731 n521 n1827 NETTRAN_DUMMY_8670 NETTRAN_DUMMY_8671 INV_X1 
XU1732 n1826 n1828 NETTRAN_DUMMY_8672 NETTRAN_DUMMY_8673 INV_X32 
XU1733 n1832 n1829 NETTRAN_DUMMY_8674 NETTRAN_DUMMY_8675 CLKBUF_X1 
XU1734 n1829 n1830 NETTRAN_DUMMY_8676 NETTRAN_DUMMY_8677 INV_X32 
XU1735 n1830 n1831 NETTRAN_DUMMY_8678 NETTRAN_DUMMY_8679 INV_X1 
XU1736 n514 n1832 NETTRAN_DUMMY_8680 NETTRAN_DUMMY_8681 INV_X1 
XU1737 n1831 n1833 NETTRAN_DUMMY_8682 NETTRAN_DUMMY_8683 INV_X32 
XU1738 n1839 n1834 NETTRAN_DUMMY_8684 NETTRAN_DUMMY_8685 INV_X1 
XU1739 n1834 n1835 NETTRAN_DUMMY_8686 NETTRAN_DUMMY_8687 INV_X32 
XU1740 n507 n1836 NETTRAN_DUMMY_8688 NETTRAN_DUMMY_8689 INV_X1 
XU1741 n1836 n1837 NETTRAN_DUMMY_8690 NETTRAN_DUMMY_8691 INV_X32 
XU1742 n1837 n1838 NETTRAN_DUMMY_8692 NETTRAN_DUMMY_8693 INV_X1 
XU1743 n1838 n1839 NETTRAN_DUMMY_8694 NETTRAN_DUMMY_8695 INV_X32 
XU1744 n1843 n1840 NETTRAN_DUMMY_8696 NETTRAN_DUMMY_8697 CLKBUF_X1 
XU1745 n1840 n1841 NETTRAN_DUMMY_8698 NETTRAN_DUMMY_8699 INV_X32 
XU1746 n1841 n1842 NETTRAN_DUMMY_8700 NETTRAN_DUMMY_8701 INV_X1 
XU1747 n500 n1843 NETTRAN_DUMMY_8702 NETTRAN_DUMMY_8703 INV_X1 
XU1748 n1842 n1844 NETTRAN_DUMMY_8704 NETTRAN_DUMMY_8705 INV_X32 
XU1749 n1848 n1845 NETTRAN_DUMMY_8706 NETTRAN_DUMMY_8707 CLKBUF_X1 
XU1750 n1845 n1846 NETTRAN_DUMMY_8708 NETTRAN_DUMMY_8709 INV_X32 
XU1751 n1846 n1847 NETTRAN_DUMMY_8710 NETTRAN_DUMMY_8711 INV_X1 
XU1752 n545 n1848 NETTRAN_DUMMY_8712 NETTRAN_DUMMY_8713 INV_X1 
XU1753 n1847 n1849 NETTRAN_DUMMY_8714 NETTRAN_DUMMY_8715 INV_X32 
XU1754 n1851 n1850 NETTRAN_DUMMY_8716 NETTRAN_DUMMY_8717 CLKBUF_X1 
XU1755 n1854 n1851 NETTRAN_DUMMY_8718 NETTRAN_DUMMY_8719 INV_X1 
XU1756 n1850 n1852 NETTRAN_DUMMY_8720 NETTRAN_DUMMY_8721 INV_X32 
XU1757 n538 n1853 NETTRAN_DUMMY_8722 NETTRAN_DUMMY_8723 INV_X1 
XU1758 n1853 n1854 NETTRAN_DUMMY_8724 NETTRAN_DUMMY_8725 INV_X32 
XU1759 n1858 n1855 NETTRAN_DUMMY_8726 NETTRAN_DUMMY_8727 CLKBUF_X1 
XU1760 n531 n1856 NETTRAN_DUMMY_8728 NETTRAN_DUMMY_8729 INV_X1 
XU1761 n1856 n1857 NETTRAN_DUMMY_8730 NETTRAN_DUMMY_8731 INV_X32 
XU1762 n1857 n1858 NETTRAN_DUMMY_8732 NETTRAN_DUMMY_8733 INV_X1 
XU1763 n1855 n1859 NETTRAN_DUMMY_8734 NETTRAN_DUMMY_8735 INV_X32 
XU1764 n1865 n1860 NETTRAN_DUMMY_8736 NETTRAN_DUMMY_8737 INV_X1 
XU1765 n1860 n1861 NETTRAN_DUMMY_8738 NETTRAN_DUMMY_8739 INV_X32 
XU1766 n1864 n1862 NETTRAN_DUMMY_8740 NETTRAN_DUMMY_8741 INV_X32 
XU1767 n1862 n1863 NETTRAN_DUMMY_8742 NETTRAN_DUMMY_8743 INV_X1 
XU1768 n524 n1864 NETTRAN_DUMMY_8744 NETTRAN_DUMMY_8745 INV_X1 
XU1769 n1863 n1865 NETTRAN_DUMMY_8746 NETTRAN_DUMMY_8747 INV_X32 
XU1770 n1867 n1866 NETTRAN_DUMMY_8748 NETTRAN_DUMMY_8749 CLKBUF_X1 
XU1771 n1870 n1867 NETTRAN_DUMMY_8750 NETTRAN_DUMMY_8751 INV_X1 
XU1772 n1866 n1868 NETTRAN_DUMMY_8752 NETTRAN_DUMMY_8753 INV_X32 
XU1773 n517 n1869 NETTRAN_DUMMY_8754 NETTRAN_DUMMY_8755 INV_X1 
XU1774 n1869 n1870 NETTRAN_DUMMY_8756 NETTRAN_DUMMY_8757 INV_X32 
XU1775 n1874 n1871 NETTRAN_DUMMY_8758 NETTRAN_DUMMY_8759 CLKBUF_X1 
XU1776 n1871 n1872 NETTRAN_DUMMY_8760 NETTRAN_DUMMY_8761 INV_X32 
XU1777 n1872 n1873 NETTRAN_DUMMY_8762 NETTRAN_DUMMY_8763 INV_X1 
XU1778 n510 n1874 NETTRAN_DUMMY_8764 NETTRAN_DUMMY_8765 INV_X1 
XU1779 n1873 n1875 NETTRAN_DUMMY_8766 NETTRAN_DUMMY_8767 INV_X32 
XU1780 n503 n1876 NETTRAN_DUMMY_8768 NETTRAN_DUMMY_8769 INV_X1 
XU1781 n1876 n1877 NETTRAN_DUMMY_8770 NETTRAN_DUMMY_8771 INV_X32 
XU1782 n1877 n1878 NETTRAN_DUMMY_8772 NETTRAN_DUMMY_8773 INV_X1 
XU1783 n723 n1879 NETTRAN_DUMMY_8774 NETTRAN_DUMMY_8775 INV_X32 
XU1784 n7 n1880 NETTRAN_DUMMY_8776 NETTRAN_DUMMY_8777 INV_X1 
XU1785 n1880 n1881 NETTRAN_DUMMY_8778 NETTRAN_DUMMY_8779 INV_X8 
XU1786 n725 n1882 NETTRAN_DUMMY_8780 NETTRAN_DUMMY_8781 INV_X32 
XU1787 n1882 n1883 NETTRAN_DUMMY_8782 NETTRAN_DUMMY_8783 INV_X1 
XU1788 n548 n1884 NETTRAN_DUMMY_8784 NETTRAN_DUMMY_8785 INV_X1 
XU1789 n1883 n1885 NETTRAN_DUMMY_8786 NETTRAN_DUMMY_8787 INV_X32 
XU1790 n52 n1886 NETTRAN_DUMMY_8788 NETTRAN_DUMMY_8789 CLKBUF_X1 
XU1791 n1888 n1887 NETTRAN_DUMMY_8790 NETTRAN_DUMMY_8791 CLKBUF_X1 
XU1792 n541 n1888 NETTRAN_DUMMY_8792 NETTRAN_DUMMY_8793 INV_X1 
XU1793 n1887 n1889 NETTRAN_DUMMY_8794 NETTRAN_DUMMY_8795 INV_X32 
XU1794 n1889 n1890 NETTRAN_DUMMY_8796 NETTRAN_DUMMY_8797 INV_X1 
XU1795 n1890 n1891 NETTRAN_DUMMY_8798 NETTRAN_DUMMY_8799 INV_X32 
XU1796 n1895 n1892 NETTRAN_DUMMY_8800 NETTRAN_DUMMY_8801 CLKBUF_X1 
XU1797 n534 n1893 NETTRAN_DUMMY_8802 NETTRAN_DUMMY_8803 INV_X1 
XU1798 n1893 n1894 NETTRAN_DUMMY_8804 NETTRAN_DUMMY_8805 INV_X32 
XU1799 n1894 n1895 NETTRAN_DUMMY_8806 NETTRAN_DUMMY_8807 INV_X1 
XU1800 n1892 n1896 NETTRAN_DUMMY_8808 NETTRAN_DUMMY_8809 INV_X32 
XU1801 n1900 n1897 NETTRAN_DUMMY_8810 NETTRAN_DUMMY_8811 CLKBUF_X1 
XU1802 n527 n1898 NETTRAN_DUMMY_8812 NETTRAN_DUMMY_8813 INV_X1 
XU1803 n1898 n1899 NETTRAN_DUMMY_8814 NETTRAN_DUMMY_8815 INV_X32 
XU1804 n1899 n1900 NETTRAN_DUMMY_8816 NETTRAN_DUMMY_8817 INV_X1 
XU1805 n1897 n1901 NETTRAN_DUMMY_8818 NETTRAN_DUMMY_8819 INV_X32 
XU1806 n1903 n1902 NETTRAN_DUMMY_8820 NETTRAN_DUMMY_8821 CLKBUF_X1 
XU1807 n1906 n1903 NETTRAN_DUMMY_8822 NETTRAN_DUMMY_8823 INV_X1 
XU1808 n1902 n1904 NETTRAN_DUMMY_8824 NETTRAN_DUMMY_8825 INV_X32 
XU1809 n520 n1905 NETTRAN_DUMMY_8826 NETTRAN_DUMMY_8827 INV_X1 
XU1810 n1905 n1906 NETTRAN_DUMMY_8828 NETTRAN_DUMMY_8829 INV_X32 
XU1811 n1908 n1907 NETTRAN_DUMMY_8830 NETTRAN_DUMMY_8831 CLKBUF_X1 
XU1812 n513 n1908 NETTRAN_DUMMY_8832 NETTRAN_DUMMY_8833 INV_X1 
XU1813 n1907 n1909 NETTRAN_DUMMY_8834 NETTRAN_DUMMY_8835 INV_X32 
XU1814 n1909 n1910 NETTRAN_DUMMY_8836 NETTRAN_DUMMY_8837 INV_X1 
XU1815 n1910 n1911 NETTRAN_DUMMY_8838 NETTRAN_DUMMY_8839 INV_X32 
XU1816 n1915 n1912 NETTRAN_DUMMY_8840 NETTRAN_DUMMY_8841 CLKBUF_X1 
XU1817 n1912 n1913 NETTRAN_DUMMY_8842 NETTRAN_DUMMY_8843 INV_X32 
XU1818 n1913 n1914 NETTRAN_DUMMY_8844 NETTRAN_DUMMY_8845 INV_X1 
XU1819 n506 n1915 NETTRAN_DUMMY_8846 NETTRAN_DUMMY_8847 INV_X1 
XU1820 n1914 n1916 NETTRAN_DUMMY_8848 NETTRAN_DUMMY_8849 INV_X32 
XU1821 n1920 n1917 NETTRAN_DUMMY_8850 NETTRAN_DUMMY_8851 CLKBUF_X1 
XU1822 n1917 n1918 NETTRAN_DUMMY_8852 NETTRAN_DUMMY_8853 INV_X32 
XU1823 n1918 n1919 NETTRAN_DUMMY_8854 NETTRAN_DUMMY_8855 INV_X1 
XU1824 n499 n1920 NETTRAN_DUMMY_8856 NETTRAN_DUMMY_8857 INV_X1 
XU1825 n1919 n1921 NETTRAN_DUMMY_8858 NETTRAN_DUMMY_8859 INV_X32 
XU1826 n1925 n1922 NETTRAN_DUMMY_8860 NETTRAN_DUMMY_8861 CLKBUF_X1 
XU1827 n1922 n1923 NETTRAN_DUMMY_8862 NETTRAN_DUMMY_8863 INV_X32 
XU1828 n1923 n1924 NETTRAN_DUMMY_8864 NETTRAN_DUMMY_8865 INV_X1 
XU1829 n496 n1925 NETTRAN_DUMMY_8866 NETTRAN_DUMMY_8867 INV_X1 
XU1830 n1924 n1926 NETTRAN_DUMMY_8868 NETTRAN_DUMMY_8869 INV_X32 
XU1831 n736 n1927 NETTRAN_DUMMY_8870 NETTRAN_DUMMY_8871 INV_X32 
XU1832 n1927 n1928 NETTRAN_DUMMY_8872 NETTRAN_DUMMY_8873 INV_X1 
XU1833 n472 n1929 NETTRAN_DUMMY_8874 NETTRAN_DUMMY_8875 INV_X1 
XU1834 n1928 n1930 NETTRAN_DUMMY_8876 NETTRAN_DUMMY_8877 INV_X32 
XU1835 n99 n1931 NETTRAN_DUMMY_8878 NETTRAN_DUMMY_8879 BUF_X1 
XU1836 n1937 n1932 NETTRAN_DUMMY_8880 NETTRAN_DUMMY_8881 INV_X1 
XU1837 n1932 n1933 NETTRAN_DUMMY_8882 NETTRAN_DUMMY_8883 INV_X32 
XU1838 n448 n1934 NETTRAN_DUMMY_8884 NETTRAN_DUMMY_8885 INV_X1 
XU1839 n1934 n1935 NETTRAN_DUMMY_8886 NETTRAN_DUMMY_8887 INV_X32 
XU1840 n1935 n1936 NETTRAN_DUMMY_8888 NETTRAN_DUMMY_8889 INV_X1 
XU1841 n1936 n1937 NETTRAN_DUMMY_8890 NETTRAN_DUMMY_8891 INV_X32 
XU1842 n1941 n1938 NETTRAN_DUMMY_8892 NETTRAN_DUMMY_8893 CLKBUF_X1 
XU1843 n482 n1939 NETTRAN_DUMMY_8894 NETTRAN_DUMMY_8895 INV_X1 
XU1844 n1939 n1940 NETTRAN_DUMMY_8896 NETTRAN_DUMMY_8897 INV_X32 
XU1845 n1940 n1941 NETTRAN_DUMMY_8898 NETTRAN_DUMMY_8899 INV_X1 
XU1846 n1938 n1942 NETTRAN_DUMMY_8900 NETTRAN_DUMMY_8901 INV_X32 
XU1847 n1946 n1943 NETTRAN_DUMMY_8902 NETTRAN_DUMMY_8903 CLKBUF_X1 
XU1848 n1943 n1944 NETTRAN_DUMMY_8904 NETTRAN_DUMMY_8905 INV_X32 
XU1849 n1944 n1945 NETTRAN_DUMMY_8906 NETTRAN_DUMMY_8907 INV_X1 
XU1850 n458 n1946 NETTRAN_DUMMY_8908 NETTRAN_DUMMY_8909 INV_X1 
XU1851 n1945 n1947 NETTRAN_DUMMY_8910 NETTRAN_DUMMY_8911 INV_X32 
XU1852 n1953 n1948 NETTRAN_DUMMY_8912 NETTRAN_DUMMY_8913 INV_X1 
XU1853 n1948 n1949 NETTRAN_DUMMY_8914 NETTRAN_DUMMY_8915 INV_X32 
XU1854 n1952 n1950 NETTRAN_DUMMY_8916 NETTRAN_DUMMY_8917 INV_X32 
XU1855 n1950 n1951 NETTRAN_DUMMY_8918 NETTRAN_DUMMY_8919 INV_X1 
XU1856 n434 n1952 NETTRAN_DUMMY_8920 NETTRAN_DUMMY_8921 INV_X1 
XU1857 n1951 n1953 NETTRAN_DUMMY_8922 NETTRAN_DUMMY_8923 INV_X32 
XU1858 n1957 n1954 NETTRAN_DUMMY_8924 NETTRAN_DUMMY_8925 CLKBUF_X1 
XU1859 n1954 n1955 NETTRAN_DUMMY_8926 NETTRAN_DUMMY_8927 INV_X32 
XU1860 n1955 n1956 NETTRAN_DUMMY_8928 NETTRAN_DUMMY_8929 INV_X1 
XU1861 n492 n1957 NETTRAN_DUMMY_8930 NETTRAN_DUMMY_8931 INV_X1 
XU1862 n1956 n1958 NETTRAN_DUMMY_8932 NETTRAN_DUMMY_8933 INV_X32 
XU1863 n1962 n1959 NETTRAN_DUMMY_8934 NETTRAN_DUMMY_8935 CLKBUF_X1 
XU1864 n1959 n1960 NETTRAN_DUMMY_8936 NETTRAN_DUMMY_8937 INV_X32 
XU1865 n1960 n1961 NETTRAN_DUMMY_8938 NETTRAN_DUMMY_8939 INV_X1 
XU1866 n468 n1962 NETTRAN_DUMMY_8940 NETTRAN_DUMMY_8941 INV_X1 
XU1867 n1961 n1963 NETTRAN_DUMMY_8942 NETTRAN_DUMMY_8943 INV_X32 
XU1868 n1967 n1964 NETTRAN_DUMMY_8944 NETTRAN_DUMMY_8945 CLKBUF_X1 
XU1869 n444 n1965 NETTRAN_DUMMY_8946 NETTRAN_DUMMY_8947 INV_X1 
XU1870 n1965 n1966 NETTRAN_DUMMY_8948 NETTRAN_DUMMY_8949 INV_X32 
XU1871 n1966 n1967 NETTRAN_DUMMY_8950 NETTRAN_DUMMY_8951 INV_X1 
XU1872 n1964 n1968 NETTRAN_DUMMY_8952 NETTRAN_DUMMY_8953 INV_X32 
XU1873 n478 n1969 NETTRAN_DUMMY_8954 NETTRAN_DUMMY_8955 INV_X1 
XU1874 n1969 n1970 NETTRAN_DUMMY_8956 NETTRAN_DUMMY_8957 INV_X32 
XU1875 n1970 n1971 NETTRAN_DUMMY_8958 NETTRAN_DUMMY_8959 INV_X1 
XU1876 n1971 n1972 NETTRAN_DUMMY_8960 NETTRAN_DUMMY_8961 INV_X32 
XU1877 n1973 n1974 NETTRAN_DUMMY_8962 NETTRAN_DUMMY_8963 INV_X1 
XU1878 n1980 n1975 NETTRAN_DUMMY_8964 NETTRAN_DUMMY_8965 INV_X1 
XU1879 n1975 n1976 NETTRAN_DUMMY_8966 NETTRAN_DUMMY_8967 INV_X32 
XU1880 n1979 n1977 NETTRAN_DUMMY_8968 NETTRAN_DUMMY_8969 INV_X32 
XU1881 n1977 n1978 NETTRAN_DUMMY_8970 NETTRAN_DUMMY_8971 INV_X1 
XU1882 n454 n1979 NETTRAN_DUMMY_8972 NETTRAN_DUMMY_8973 INV_X1 
XU1883 n1978 n1980 NETTRAN_DUMMY_8974 NETTRAN_DUMMY_8975 INV_X32 
XU1884 n1984 n1981 NETTRAN_DUMMY_8976 NETTRAN_DUMMY_8977 CLKBUF_X1 
XU1885 n1981 n1982 NETTRAN_DUMMY_8978 NETTRAN_DUMMY_8979 INV_X32 
XU1886 n1982 n1983 NETTRAN_DUMMY_8980 NETTRAN_DUMMY_8981 INV_X1 
XU1887 n493 n1984 NETTRAN_DUMMY_8982 NETTRAN_DUMMY_8983 INV_X1 
XU1888 n1983 n1985 NETTRAN_DUMMY_8984 NETTRAN_DUMMY_8985 INV_X32 
XU1889 n1987 n1986 NETTRAN_DUMMY_8986 NETTRAN_DUMMY_8987 CLKBUF_X1 
XU1890 n469 n1987 NETTRAN_DUMMY_8988 NETTRAN_DUMMY_8989 INV_X1 
XU1891 n1986 n1988 NETTRAN_DUMMY_8990 NETTRAN_DUMMY_8991 INV_X32 
XU1892 n1988 n1989 NETTRAN_DUMMY_8992 NETTRAN_DUMMY_8993 INV_X1 
XU1893 n1989 n1990 NETTRAN_DUMMY_8994 NETTRAN_DUMMY_8995 INV_X32 
XU1894 n1994 n1991 NETTRAN_DUMMY_8996 NETTRAN_DUMMY_8997 CLKBUF_X1 
XU1895 n1991 n1992 NETTRAN_DUMMY_8998 NETTRAN_DUMMY_8999 INV_X32 
XU1896 n1992 n1993 NETTRAN_DUMMY_9000 NETTRAN_DUMMY_9001 INV_X1 
XU1897 n445 n1994 NETTRAN_DUMMY_9002 NETTRAN_DUMMY_9003 INV_X1 
XU1898 n1993 n1995 NETTRAN_DUMMY_9004 NETTRAN_DUMMY_9005 INV_X32 
XU1899 n1999 n1996 NETTRAN_DUMMY_9006 NETTRAN_DUMMY_9007 INV_X1 
XU1900 n1996 n1997 NETTRAN_DUMMY_9008 NETTRAN_DUMMY_9009 INV_X32 
XU1901 n479 n1998 NETTRAN_DUMMY_9010 NETTRAN_DUMMY_9011 INV_X1 
XU1902 n1998 n1999 NETTRAN_DUMMY_9012 NETTRAN_DUMMY_9013 INV_X32 
XU1903 n106 n2000 NETTRAN_DUMMY_9014 NETTRAN_DUMMY_9015 INV_X32 
XU1904 n2000 n2001 NETTRAN_DUMMY_9016 NETTRAN_DUMMY_9017 INV_X1 
XU1905 n2005 n2002 NETTRAN_DUMMY_9018 NETTRAN_DUMMY_9019 INV_X32 
XU1906 n2002 n2003 NETTRAN_DUMMY_9020 NETTRAN_DUMMY_9021 INV_X1 
XU1907 n2006 n2004 NETTRAN_DUMMY_9022 NETTRAN_DUMMY_9023 INV_X32 
XU1908 n2004 n2005 NETTRAN_DUMMY_9024 NETTRAN_DUMMY_9025 INV_X1 
XU1909 n455 n2006 NETTRAN_DUMMY_9026 NETTRAN_DUMMY_9027 INV_X1 
XU1910 n2003 n2007 NETTRAN_DUMMY_9028 NETTRAN_DUMMY_9029 INV_X32 
XU1911 n2011 n2008 NETTRAN_DUMMY_9030 NETTRAN_DUMMY_9031 CLKBUF_X1 
XU1912 n2008 n2009 NETTRAN_DUMMY_9032 NETTRAN_DUMMY_9033 INV_X32 
XU1913 n2009 n2010 NETTRAN_DUMMY_9034 NETTRAN_DUMMY_9035 INV_X1 
XU1914 n494 n2011 NETTRAN_DUMMY_9036 NETTRAN_DUMMY_9037 INV_X1 
XU1915 n2010 n2012 NETTRAN_DUMMY_9038 NETTRAN_DUMMY_9039 INV_X32 
XU1916 n2025 n2013 NETTRAN_DUMMY_9040 NETTRAN_DUMMY_9041 CLKBUF_X1 
XU1917 n2015 n2014 NETTRAN_DUMMY_9042 NETTRAN_DUMMY_9043 CLKBUF_X1 
XU1918 n2013 n2015 NETTRAN_DUMMY_9044 NETTRAN_DUMMY_9045 INV_X32 
XU1919 n2014 data_out[0] NETTRAN_DUMMY_9046 NETTRAN_DUMMY_9047 INV_X32 
XU1920 n2026 n2017 NETTRAN_DUMMY_9048 NETTRAN_DUMMY_9049 CLKBUF_X1 
XU1921 n2017 n2018 NETTRAN_DUMMY_9050 NETTRAN_DUMMY_9051 INV_X32 
XU1922 n2018 data_out[6] NETTRAN_DUMMY_9052 NETTRAN_DUMMY_9053 INV_X1 
XU1923 n2024 n2020 NETTRAN_DUMMY_9054 NETTRAN_DUMMY_9055 CLKBUF_X1 
XU1924 n2022 n2021 NETTRAN_DUMMY_9056 NETTRAN_DUMMY_9057 CLKBUF_X1 
XU1925 n2020 n2022 NETTRAN_DUMMY_9058 NETTRAN_DUMMY_9059 INV_X32 
XU1926 n2021 data_out[14] NETTRAN_DUMMY_9060 NETTRAN_DUMMY_9061 INV_X32 
XU722 n811 n812 NETTRAN_DUMMY_9062 NETTRAN_DUMMY_9063 INV_X2 
XU1927 n812 n2027 NETTRAN_DUMMY_9064 NETTRAN_DUMMY_9065 BUF_X1 
XU1928 n1071 n2028 NETTRAN_DUMMY_9066 NETTRAN_DUMMY_9067 BUF_X1 
XU1929 n830 n2029 NETTRAN_DUMMY_9068 NETTRAN_DUMMY_9069 BUF_X1 
XU1930 n1045 n2030 NETTRAN_DUMMY_9070 NETTRAN_DUMMY_9071 BUF_X1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW01_add_1 CI CO SUM[31] SUM[30] SUM[29] SUM[28] SUM[27] 
+ SUM[26] SUM[25] SUM[24] SUM[23] SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] SUM[17] 
+ SUM[16] SUM[15] SUM[14] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] B[23] 
+ B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] 
+ B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[31] A[30] A[29] A[28] A[27] 
+ A[26] A[25] A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] 
+ A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU7 n30 n3 NETTRAN_DUMMY_9072 NETTRAN_DUMMY_9073 INV_X1 
XU6 n38 n5 NETTRAN_DUMMY_9074 NETTRAN_DUMMY_9075 INV_X1 
XU5 n46 n7 NETTRAN_DUMMY_9076 NETTRAN_DUMMY_9077 INV_X1 
XU4 n54 n9 NETTRAN_DUMMY_9078 NETTRAN_DUMMY_9079 INV_X1 
XU3 n62 n11 NETTRAN_DUMMY_9080 NETTRAN_DUMMY_9081 INV_X1 
XU2 n70 n13 NETTRAN_DUMMY_9082 NETTRAN_DUMMY_9083 INV_X1 
XU100 B[15] A[15] n80 NETTRAN_DUMMY_9084 NETTRAN_DUMMY_9085 NOR2_X1 
XU99 B[15] A[15] n82 NETTRAN_DUMMY_9086 NETTRAN_DUMMY_9087 NAND2_X1 
XU98 n16 n82 n83 NETTRAN_DUMMY_9088 NETTRAN_DUMMY_9089 NAND2_X1 
XU97 n81 n83 n155 NETTRAN_DUMMY_9090 NETTRAN_DUMMY_9091 XOR2_X1 
XU96 n82 n80 n81 n76 NETTRAN_DUMMY_9092 NETTRAN_DUMMY_9093 OAI21_X1 
XU95 B[16] A[16] n77 NETTRAN_DUMMY_9094 NETTRAN_DUMMY_9095 AND2_X1 
XU94 B[16] A[16] n78 NETTRAN_DUMMY_9096 NETTRAN_DUMMY_9097 NOR2_X1 
XU93 n77 n78 n79 NETTRAN_DUMMY_9098 NETTRAN_DUMMY_9099 NOR2_X1 
XU92 n76 n79 n147 NETTRAN_DUMMY_9100 NETTRAN_DUMMY_9101 XOR2_X1 
XU91 B[17] A[17] n72 NETTRAN_DUMMY_9102 NETTRAN_DUMMY_9103 NOR2_X1 
XU90 B[17] A[17] n74 NETTRAN_DUMMY_9104 NETTRAN_DUMMY_9105 NAND2_X1 
XU89 n14 n74 n75 NETTRAN_DUMMY_9106 NETTRAN_DUMMY_9107 NAND2_X1 
XU88 n77 n15 n76 n73 NETTRAN_DUMMY_9108 NETTRAN_DUMMY_9109 AOI21_X1 
XU87 n75 n73 n148 NETTRAN_DUMMY_9110 NETTRAN_DUMMY_9111 XOR2_X1 
XU86 n74 n72 n73 n68 NETTRAN_DUMMY_9112 NETTRAN_DUMMY_9113 OAI21_X1 
XU85 B[18] A[18] n69 NETTRAN_DUMMY_9114 NETTRAN_DUMMY_9115 AND2_X1 
XU84 B[18] A[18] n70 NETTRAN_DUMMY_9116 NETTRAN_DUMMY_9117 NOR2_X1 
XU83 n69 n70 n71 NETTRAN_DUMMY_9118 NETTRAN_DUMMY_9119 NOR2_X1 
XU82 n68 n71 n149 NETTRAN_DUMMY_9120 NETTRAN_DUMMY_9121 XOR2_X1 
XU81 B[19] A[19] n64 NETTRAN_DUMMY_9122 NETTRAN_DUMMY_9123 NOR2_X1 
XU80 B[19] A[19] n66 NETTRAN_DUMMY_9124 NETTRAN_DUMMY_9125 NAND2_X1 
XU79 n12 n66 n67 NETTRAN_DUMMY_9126 NETTRAN_DUMMY_9127 NAND2_X1 
XU78 n69 n13 n68 n65 NETTRAN_DUMMY_9128 NETTRAN_DUMMY_9129 AOI21_X1 
XU77 n67 n65 n150 NETTRAN_DUMMY_9130 NETTRAN_DUMMY_9131 XOR2_X1 
XU76 n66 n64 n65 n60 NETTRAN_DUMMY_9132 NETTRAN_DUMMY_9133 OAI21_X1 
XU75 B[20] A[20] n61 NETTRAN_DUMMY_9134 NETTRAN_DUMMY_9135 AND2_X1 
XU74 B[20] A[20] n62 NETTRAN_DUMMY_9136 NETTRAN_DUMMY_9137 NOR2_X1 
XU73 n61 n62 n63 NETTRAN_DUMMY_9138 NETTRAN_DUMMY_9139 NOR2_X1 
XU72 n60 n63 n151 NETTRAN_DUMMY_9140 NETTRAN_DUMMY_9141 XOR2_X1 
XU71 B[21] A[21] n56 NETTRAN_DUMMY_9142 NETTRAN_DUMMY_9143 NOR2_X1 
XU70 B[21] A[21] n58 NETTRAN_DUMMY_9144 NETTRAN_DUMMY_9145 NAND2_X1 
XU69 n10 n58 n59 NETTRAN_DUMMY_9146 NETTRAN_DUMMY_9147 NAND2_X1 
XU68 n61 n11 n60 n57 NETTRAN_DUMMY_9148 NETTRAN_DUMMY_9149 AOI21_X1 
XU67 n59 n57 n152 NETTRAN_DUMMY_9150 NETTRAN_DUMMY_9151 XOR2_X1 
XU66 n58 n56 n57 n52 NETTRAN_DUMMY_9152 NETTRAN_DUMMY_9153 OAI21_X1 
XU65 B[22] A[22] n53 NETTRAN_DUMMY_9154 NETTRAN_DUMMY_9155 AND2_X1 
XU64 B[22] A[22] n54 NETTRAN_DUMMY_9156 NETTRAN_DUMMY_9157 NOR2_X1 
XU63 n53 n54 n55 NETTRAN_DUMMY_9158 NETTRAN_DUMMY_9159 NOR2_X1 
XU62 n52 n55 n153 NETTRAN_DUMMY_9160 NETTRAN_DUMMY_9161 XOR2_X1 
XU61 B[23] A[23] n48 NETTRAN_DUMMY_9162 NETTRAN_DUMMY_9163 NOR2_X1 
XU60 B[23] A[23] n50 NETTRAN_DUMMY_9164 NETTRAN_DUMMY_9165 NAND2_X1 
XU59 n8 n85 n51 NETTRAN_DUMMY_9166 NETTRAN_DUMMY_9167 NAND2_X1 
XU58 n53 n9 n52 n49 NETTRAN_DUMMY_9168 NETTRAN_DUMMY_9169 AOI21_X1 
XU57 n51 n49 n154 NETTRAN_DUMMY_9170 NETTRAN_DUMMY_9171 XOR2_X1 
XU56 n85 n48 n49 n44 NETTRAN_DUMMY_9172 NETTRAN_DUMMY_9173 OAI21_X1 
XU55 B[24] A[24] n45 NETTRAN_DUMMY_9174 NETTRAN_DUMMY_9175 AND2_X1 
XU54 B[24] A[24] n46 NETTRAN_DUMMY_9176 NETTRAN_DUMMY_9177 NOR2_X1 
XU53 n45 n46 n47 NETTRAN_DUMMY_9178 NETTRAN_DUMMY_9179 NOR2_X1 
XU52 n44 n47 n139 NETTRAN_DUMMY_9180 NETTRAN_DUMMY_9181 XOR2_X1 
XU51 B[25] A[25] n40 NETTRAN_DUMMY_9182 NETTRAN_DUMMY_9183 NOR2_X1 
XU50 B[25] A[25] n42 NETTRAN_DUMMY_9184 NETTRAN_DUMMY_9185 NAND2_X1 
XU49 n6 n42 n43 NETTRAN_DUMMY_9186 NETTRAN_DUMMY_9187 NAND2_X1 
XU48 n45 n7 n44 n41 NETTRAN_DUMMY_9188 NETTRAN_DUMMY_9189 AOI21_X1 
XU47 n43 n41 n140 NETTRAN_DUMMY_9190 NETTRAN_DUMMY_9191 XOR2_X1 
XU46 n42 n40 n41 n36 NETTRAN_DUMMY_9192 NETTRAN_DUMMY_9193 OAI21_X1 
XU45 B[26] A[26] n37 NETTRAN_DUMMY_9194 NETTRAN_DUMMY_9195 AND2_X1 
XU44 B[26] A[26] n38 NETTRAN_DUMMY_9196 NETTRAN_DUMMY_9197 NOR2_X1 
XU43 n37 n38 n39 NETTRAN_DUMMY_9198 NETTRAN_DUMMY_9199 NOR2_X1 
XU42 n36 n39 n141 NETTRAN_DUMMY_9200 NETTRAN_DUMMY_9201 XOR2_X1 
XU41 B[27] A[27] n32 NETTRAN_DUMMY_9202 NETTRAN_DUMMY_9203 NOR2_X1 
XU40 B[27] A[27] n34 NETTRAN_DUMMY_9204 NETTRAN_DUMMY_9205 NAND2_X1 
XU39 n4 n34 n35 NETTRAN_DUMMY_9206 NETTRAN_DUMMY_9207 NAND2_X1 
XU38 n37 n5 n36 n33 NETTRAN_DUMMY_9208 NETTRAN_DUMMY_9209 AOI21_X1 
XU37 n35 n33 n142 NETTRAN_DUMMY_9210 NETTRAN_DUMMY_9211 XOR2_X1 
XU36 n34 n32 n33 n28 NETTRAN_DUMMY_9212 NETTRAN_DUMMY_9213 OAI21_X1 
XU35 B[28] A[28] n29 NETTRAN_DUMMY_9214 NETTRAN_DUMMY_9215 AND2_X1 
XU34 B[28] A[28] n30 NETTRAN_DUMMY_9216 NETTRAN_DUMMY_9217 NOR2_X1 
XU33 n29 n30 n31 NETTRAN_DUMMY_9218 NETTRAN_DUMMY_9219 NOR2_X1 
XU32 n28 n31 n143 NETTRAN_DUMMY_9220 NETTRAN_DUMMY_9221 XOR2_X1 
XU31 B[29] A[29] n24 NETTRAN_DUMMY_9222 NETTRAN_DUMMY_9223 NOR2_X1 
XU30 B[29] A[29] n26 NETTRAN_DUMMY_9224 NETTRAN_DUMMY_9225 NAND2_X1 
XU29 n2 n26 n27 NETTRAN_DUMMY_9226 NETTRAN_DUMMY_9227 NAND2_X1 
XU28 n29 n3 n28 n25 NETTRAN_DUMMY_9228 NETTRAN_DUMMY_9229 AOI21_X1 
XU27 n27 n25 n144 NETTRAN_DUMMY_9230 NETTRAN_DUMMY_9231 XOR2_X1 
XU26 n26 n24 n25 n20 NETTRAN_DUMMY_9232 NETTRAN_DUMMY_9233 OAI21_X1 
XU25 B[30] A[30] n21 NETTRAN_DUMMY_9234 NETTRAN_DUMMY_9235 AND2_X1 
XU24 B[30] A[30] n22 NETTRAN_DUMMY_9236 NETTRAN_DUMMY_9237 NOR2_X1 
XU23 n21 n22 n23 NETTRAN_DUMMY_9238 NETTRAN_DUMMY_9239 NOR2_X1 
XU22 n20 n23 n145 NETTRAN_DUMMY_9240 NETTRAN_DUMMY_9241 XOR2_X1 
XU21 B[31] A[31] n18 NETTRAN_DUMMY_9242 NETTRAN_DUMMY_9243 XNOR2_X1 
XU20 n21 n20 n1 n19 NETTRAN_DUMMY_9244 NETTRAN_DUMMY_9245 AOI21_X1 
XU19 n18 n19 n146 NETTRAN_DUMMY_9246 NETTRAN_DUMMY_9247 XOR2_X1 
XU18 n126 SUM[14] NETTRAN_DUMMY_9248 NETTRAN_DUMMY_9249 INV_X1 
XU17 n80 n16 NETTRAN_DUMMY_9250 NETTRAN_DUMMY_9251 INV_X1 
XU16 n78 n15 NETTRAN_DUMMY_9252 NETTRAN_DUMMY_9253 INV_X1 
XU15 n22 n1 NETTRAN_DUMMY_9254 NETTRAN_DUMMY_9255 INV_X1 
XU14 n40 n6 NETTRAN_DUMMY_9256 NETTRAN_DUMMY_9257 INV_X1 
XU13 n48 n8 NETTRAN_DUMMY_9258 NETTRAN_DUMMY_9259 INV_X1 
XU12 n56 n10 NETTRAN_DUMMY_9260 NETTRAN_DUMMY_9261 INV_X1 
XU11 n64 n12 NETTRAN_DUMMY_9262 NETTRAN_DUMMY_9263 INV_X1 
XU10 n72 n14 NETTRAN_DUMMY_9264 NETTRAN_DUMMY_9265 INV_X1 
XU9 n24 n2 NETTRAN_DUMMY_9266 NETTRAN_DUMMY_9267 INV_X1 
XU8 n32 n4 NETTRAN_DUMMY_9268 NETTRAN_DUMMY_9269 INV_X1 
XU102 B[14] A[14] n81 NETTRAN_DUMMY_9270 NETTRAN_DUMMY_9271 NAND2_X1 
XU101 n81 B[14] A[14] n84 NETTRAN_DUMMY_9272 NETTRAN_DUMMY_9273 OAI21_X1 
XU1 n91 SUM[26] NETTRAN_DUMMY_9274 NETTRAN_DUMMY_9275 BUF_X1 
XU103 n50 n85 NETTRAN_DUMMY_9276 NETTRAN_DUMMY_9277 BUF_X1 
XU104 n107 SUM[20] NETTRAN_DUMMY_9278 NETTRAN_DUMMY_9279 BUF_X1 
XU105 n143 n137 NETTRAN_DUMMY_9280 NETTRAN_DUMMY_9281 INV_X2 
XU106 n145 n131 NETTRAN_DUMMY_9282 NETTRAN_DUMMY_9283 INV_X4 
XU107 n144 n134 NETTRAN_DUMMY_9284 NETTRAN_DUMMY_9285 INV_X4 
XU108 n153 n102 NETTRAN_DUMMY_9286 NETTRAN_DUMMY_9287 INV_X1 
XU109 n154 n99 NETTRAN_DUMMY_9288 NETTRAN_DUMMY_9289 INV_X1 
XU110 n89 n87 NETTRAN_DUMMY_9290 NETTRAN_DUMMY_9291 INV_X1 
XU111 n87 SUM[27] NETTRAN_DUMMY_9292 NETTRAN_DUMMY_9293 INV_X8 
XU112 n142 n89 NETTRAN_DUMMY_9294 NETTRAN_DUMMY_9295 BUF_X32 
XU113 n92 n90 NETTRAN_DUMMY_9296 NETTRAN_DUMMY_9297 INV_X1 
XU114 n90 n91 NETTRAN_DUMMY_9298 NETTRAN_DUMMY_9299 INV_X4 
XU115 n141 n92 NETTRAN_DUMMY_9300 NETTRAN_DUMMY_9301 BUF_X32 
XU116 n95 n93 NETTRAN_DUMMY_9302 NETTRAN_DUMMY_9303 INV_X1 
XU117 n93 SUM[25] NETTRAN_DUMMY_9304 NETTRAN_DUMMY_9305 INV_X8 
XU118 n140 n95 NETTRAN_DUMMY_9306 NETTRAN_DUMMY_9307 BUF_X32 
XU119 n97 SUM[24] NETTRAN_DUMMY_9308 NETTRAN_DUMMY_9309 BUF_X1 
XU120 n139 n97 NETTRAN_DUMMY_9310 NETTRAN_DUMMY_9311 BUF_X32 
XU121 n100 SUM[23] NETTRAN_DUMMY_9312 NETTRAN_DUMMY_9313 BUF_X1 
XU122 n99 n100 NETTRAN_DUMMY_9314 NETTRAN_DUMMY_9315 INV_X32 
XU123 n103 SUM[22] NETTRAN_DUMMY_9316 NETTRAN_DUMMY_9317 BUF_X1 
XU124 n102 n103 NETTRAN_DUMMY_9318 NETTRAN_DUMMY_9319 INV_X32 
XU125 n106 n104 NETTRAN_DUMMY_9320 NETTRAN_DUMMY_9321 INV_X1 
XU126 n104 SUM[21] NETTRAN_DUMMY_9322 NETTRAN_DUMMY_9323 INV_X8 
XU127 n152 n106 NETTRAN_DUMMY_9324 NETTRAN_DUMMY_9325 BUF_X32 
XU128 n108 n107 NETTRAN_DUMMY_9326 NETTRAN_DUMMY_9327 CLKBUF_X1 
XU129 n151 n108 NETTRAN_DUMMY_9328 NETTRAN_DUMMY_9329 BUF_X32 
XU130 n111 n109 NETTRAN_DUMMY_9330 NETTRAN_DUMMY_9331 INV_X1 
XU131 n109 SUM[19] NETTRAN_DUMMY_9332 NETTRAN_DUMMY_9333 INV_X8 
XU132 n150 n111 NETTRAN_DUMMY_9334 NETTRAN_DUMMY_9335 BUF_X32 
XU133 n114 n112 NETTRAN_DUMMY_9336 NETTRAN_DUMMY_9337 INV_X1 
XU134 n112 SUM[18] NETTRAN_DUMMY_9338 NETTRAN_DUMMY_9339 INV_X8 
XU135 n149 n114 NETTRAN_DUMMY_9340 NETTRAN_DUMMY_9341 BUF_X32 
XU136 n117 n115 NETTRAN_DUMMY_9342 NETTRAN_DUMMY_9343 INV_X1 
XU137 n115 SUM[17] NETTRAN_DUMMY_9344 NETTRAN_DUMMY_9345 INV_X8 
XU138 n148 n117 NETTRAN_DUMMY_9346 NETTRAN_DUMMY_9347 BUF_X32 
XU139 n120 SUM[16] NETTRAN_DUMMY_9348 NETTRAN_DUMMY_9349 BUF_X1 
XU140 n147 n119 NETTRAN_DUMMY_9350 NETTRAN_DUMMY_9351 INV_X1 
XU141 n119 n120 NETTRAN_DUMMY_9352 NETTRAN_DUMMY_9353 INV_X32 
XU142 n123 SUM[15] NETTRAN_DUMMY_9354 NETTRAN_DUMMY_9355 BUF_X1 
XU143 n155 n122 NETTRAN_DUMMY_9356 NETTRAN_DUMMY_9357 INV_X1 
XU144 n122 n123 NETTRAN_DUMMY_9358 NETTRAN_DUMMY_9359 INV_X32 
XU145 n125 n124 NETTRAN_DUMMY_9360 NETTRAN_DUMMY_9361 CLKBUF_X1 
XU146 n84 n125 NETTRAN_DUMMY_9362 NETTRAN_DUMMY_9363 INV_X1 
XU147 n124 n126 NETTRAN_DUMMY_9364 NETTRAN_DUMMY_9365 INV_X32 
XU148 n128 n127 NETTRAN_DUMMY_9366 NETTRAN_DUMMY_9367 CLKBUF_X1 
XU149 n146 n128 NETTRAN_DUMMY_9368 NETTRAN_DUMMY_9369 INV_X1 
XU150 n127 SUM[31] NETTRAN_DUMMY_9370 NETTRAN_DUMMY_9371 INV_X32 
XU151 n131 n130 NETTRAN_DUMMY_9372 NETTRAN_DUMMY_9373 BUF_X1 
XU152 n130 SUM[30] NETTRAN_DUMMY_9374 NETTRAN_DUMMY_9375 INV_X32 
XU153 n134 n133 NETTRAN_DUMMY_9376 NETTRAN_DUMMY_9377 BUF_X1 
XU154 n133 SUM[29] NETTRAN_DUMMY_9378 NETTRAN_DUMMY_9379 INV_X32 
XU155 n137 n136 NETTRAN_DUMMY_9380 NETTRAN_DUMMY_9381 BUF_X1 
XU156 n136 SUM[28] NETTRAN_DUMMY_9382 NETTRAN_DUMMY_9383 INV_X32 
.ENDS

.SUBCKT gng_smul_16_18_DW01_add_0 CI CO SUM[31] SUM[30] SUM[29] SUM[28] SUM[27] SUM[26] 
+ SUM[25] SUM[24] SUM[23] SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] SUM[17] SUM[16] 
+ SUM[15] SUM[14] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] B[23] B[22] B[21] 
+ B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] 
+ B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[31] A[30] A[29] A[28] A[27] A[26] A[25] A[24] 
+ A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] A[13] A[12] A[11] 
+ A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU44 B[26] A[26] n38 NETTRAN_DUMMY_9384 NETTRAN_DUMMY_9385 NOR2_X1 
XU43 n37 n38 n39 NETTRAN_DUMMY_9386 NETTRAN_DUMMY_9387 NOR2_X1 
XU42 n36 n39 n129 NETTRAN_DUMMY_9388 NETTRAN_DUMMY_9389 XOR2_X1 
XU41 B[27] A[27] n32 NETTRAN_DUMMY_9390 NETTRAN_DUMMY_9391 NOR2_X1 
XU40 B[27] A[27] n34 NETTRAN_DUMMY_9392 NETTRAN_DUMMY_9393 NAND2_X1 
XU39 n4 n34 n35 NETTRAN_DUMMY_9394 NETTRAN_DUMMY_9395 NAND2_X1 
XU38 n37 n5 n36 n33 NETTRAN_DUMMY_9396 NETTRAN_DUMMY_9397 AOI21_X1 
XU37 n35 n33 n130 NETTRAN_DUMMY_9398 NETTRAN_DUMMY_9399 XOR2_X1 
XU36 n34 n32 n33 n28 NETTRAN_DUMMY_9400 NETTRAN_DUMMY_9401 OAI21_X1 
XU35 B[28] A[28] n29 NETTRAN_DUMMY_9402 NETTRAN_DUMMY_9403 AND2_X1 
XU34 B[28] A[28] n30 NETTRAN_DUMMY_9404 NETTRAN_DUMMY_9405 NOR2_X1 
XU33 n29 n30 n31 NETTRAN_DUMMY_9406 NETTRAN_DUMMY_9407 NOR2_X1 
XU32 n28 n31 n131 NETTRAN_DUMMY_9408 NETTRAN_DUMMY_9409 XOR2_X1 
XU31 B[29] A[29] n24 NETTRAN_DUMMY_9410 NETTRAN_DUMMY_9411 NOR2_X1 
XU30 B[29] A[29] n26 NETTRAN_DUMMY_9412 NETTRAN_DUMMY_9413 NAND2_X1 
XU29 n2 n26 n27 NETTRAN_DUMMY_9414 NETTRAN_DUMMY_9415 NAND2_X1 
XU28 n29 n3 n28 n25 NETTRAN_DUMMY_9416 NETTRAN_DUMMY_9417 AOI21_X1 
XU27 n27 n25 n132 NETTRAN_DUMMY_9418 NETTRAN_DUMMY_9419 XOR2_X1 
XU26 n26 n24 n25 n20 NETTRAN_DUMMY_9420 NETTRAN_DUMMY_9421 OAI21_X1 
XU25 B[30] A[30] n21 NETTRAN_DUMMY_9422 NETTRAN_DUMMY_9423 AND2_X1 
XU24 B[30] A[30] n22 NETTRAN_DUMMY_9424 NETTRAN_DUMMY_9425 NOR2_X1 
XU23 n21 n22 n23 NETTRAN_DUMMY_9426 NETTRAN_DUMMY_9427 NOR2_X1 
XU22 n20 n23 n133 NETTRAN_DUMMY_9428 NETTRAN_DUMMY_9429 XOR2_X1 
XU21 B[31] A[31] n18 NETTRAN_DUMMY_9430 NETTRAN_DUMMY_9431 XNOR2_X1 
XU20 n21 n20 n1 n19 NETTRAN_DUMMY_9432 NETTRAN_DUMMY_9433 AOI21_X1 
XU19 n18 n19 SUM[31] NETTRAN_DUMMY_9434 NETTRAN_DUMMY_9435 XOR2_X1 
XU18 n84 SUM[14] NETTRAN_DUMMY_9436 NETTRAN_DUMMY_9437 INV_X1 
XU17 n80 n16 NETTRAN_DUMMY_9438 NETTRAN_DUMMY_9439 INV_X1 
XU16 n78 n15 NETTRAN_DUMMY_9440 NETTRAN_DUMMY_9441 INV_X1 
XU15 n22 n1 NETTRAN_DUMMY_9442 NETTRAN_DUMMY_9443 INV_X1 
XU14 n40 n6 NETTRAN_DUMMY_9444 NETTRAN_DUMMY_9445 INV_X1 
XU13 n48 n8 NETTRAN_DUMMY_9446 NETTRAN_DUMMY_9447 INV_X1 
XU12 n56 n10 NETTRAN_DUMMY_9448 NETTRAN_DUMMY_9449 INV_X1 
XU11 n64 n12 NETTRAN_DUMMY_9450 NETTRAN_DUMMY_9451 INV_X1 
XU10 n72 n14 NETTRAN_DUMMY_9452 NETTRAN_DUMMY_9453 INV_X1 
XU9 n24 n2 NETTRAN_DUMMY_9454 NETTRAN_DUMMY_9455 INV_X1 
XU8 n32 n4 NETTRAN_DUMMY_9456 NETTRAN_DUMMY_9457 INV_X1 
XU7 n30 n3 NETTRAN_DUMMY_9458 NETTRAN_DUMMY_9459 INV_X1 
XU6 n38 n5 NETTRAN_DUMMY_9460 NETTRAN_DUMMY_9461 INV_X1 
XU5 n46 n7 NETTRAN_DUMMY_9462 NETTRAN_DUMMY_9463 INV_X1 
XU4 n54 n9 NETTRAN_DUMMY_9464 NETTRAN_DUMMY_9465 INV_X1 
XU3 n62 n11 NETTRAN_DUMMY_9466 NETTRAN_DUMMY_9467 INV_X1 
XU2 n70 n13 NETTRAN_DUMMY_9468 NETTRAN_DUMMY_9469 INV_X1 
XU102 B[14] A[14] n81 NETTRAN_DUMMY_9470 NETTRAN_DUMMY_9471 NAND2_X1 
XU101 n81 B[14] A[14] n84 NETTRAN_DUMMY_9472 NETTRAN_DUMMY_9473 OAI21_X1 
XU100 B[15] A[15] n80 NETTRAN_DUMMY_9474 NETTRAN_DUMMY_9475 NOR2_X1 
XU99 B[15] A[15] n82 NETTRAN_DUMMY_9476 NETTRAN_DUMMY_9477 NAND2_X1 
XU98 n16 n82 n83 NETTRAN_DUMMY_9478 NETTRAN_DUMMY_9479 NAND2_X1 
XU97 n81 n83 SUM[15] NETTRAN_DUMMY_9480 NETTRAN_DUMMY_9481 XOR2_X1 
XU96 n82 n80 n81 n76 NETTRAN_DUMMY_9482 NETTRAN_DUMMY_9483 OAI21_X1 
XU95 B[16] A[16] n77 NETTRAN_DUMMY_9484 NETTRAN_DUMMY_9485 AND2_X1 
XU94 B[16] A[16] n78 NETTRAN_DUMMY_9486 NETTRAN_DUMMY_9487 NOR2_X1 
XU93 n77 n78 n79 NETTRAN_DUMMY_9488 NETTRAN_DUMMY_9489 NOR2_X1 
XU92 n76 n79 SUM[16] NETTRAN_DUMMY_9490 NETTRAN_DUMMY_9491 XOR2_X1 
XU91 B[17] A[17] n72 NETTRAN_DUMMY_9492 NETTRAN_DUMMY_9493 NOR2_X1 
XU90 B[17] A[17] n74 NETTRAN_DUMMY_9494 NETTRAN_DUMMY_9495 NAND2_X1 
XU89 n14 n74 n75 NETTRAN_DUMMY_9496 NETTRAN_DUMMY_9497 NAND2_X1 
XU88 n77 n15 n76 n73 NETTRAN_DUMMY_9498 NETTRAN_DUMMY_9499 AOI21_X1 
XU87 n75 n73 n134 NETTRAN_DUMMY_9500 NETTRAN_DUMMY_9501 XOR2_X1 
XU86 n74 n72 n73 n68 NETTRAN_DUMMY_9502 NETTRAN_DUMMY_9503 OAI21_X1 
XU85 B[18] A[18] n69 NETTRAN_DUMMY_9504 NETTRAN_DUMMY_9505 AND2_X1 
XU84 B[18] A[18] n70 NETTRAN_DUMMY_9506 NETTRAN_DUMMY_9507 NOR2_X1 
XU83 n69 n70 n71 NETTRAN_DUMMY_9508 NETTRAN_DUMMY_9509 NOR2_X1 
XU82 n68 n71 n135 NETTRAN_DUMMY_9510 NETTRAN_DUMMY_9511 XOR2_X1 
XU81 B[19] A[19] n64 NETTRAN_DUMMY_9512 NETTRAN_DUMMY_9513 NOR2_X1 
XU80 B[19] A[19] n66 NETTRAN_DUMMY_9514 NETTRAN_DUMMY_9515 NAND2_X1 
XU79 n12 n66 n67 NETTRAN_DUMMY_9516 NETTRAN_DUMMY_9517 NAND2_X1 
XU78 n69 n13 n68 n65 NETTRAN_DUMMY_9518 NETTRAN_DUMMY_9519 AOI21_X1 
XU77 n67 n65 n136 NETTRAN_DUMMY_9520 NETTRAN_DUMMY_9521 XOR2_X1 
XU76 n66 n64 n65 n60 NETTRAN_DUMMY_9522 NETTRAN_DUMMY_9523 OAI21_X1 
XU75 B[20] A[20] n61 NETTRAN_DUMMY_9524 NETTRAN_DUMMY_9525 AND2_X1 
XU74 B[20] A[20] n62 NETTRAN_DUMMY_9526 NETTRAN_DUMMY_9527 NOR2_X1 
XU73 n61 n62 n63 NETTRAN_DUMMY_9528 NETTRAN_DUMMY_9529 NOR2_X1 
XU72 n60 n63 n137 NETTRAN_DUMMY_9530 NETTRAN_DUMMY_9531 XOR2_X1 
XU71 B[21] A[21] n56 NETTRAN_DUMMY_9532 NETTRAN_DUMMY_9533 NOR2_X1 
XU70 B[21] A[21] n58 NETTRAN_DUMMY_9534 NETTRAN_DUMMY_9535 NAND2_X1 
XU69 n10 n58 n59 NETTRAN_DUMMY_9536 NETTRAN_DUMMY_9537 NAND2_X1 
XU68 n61 n11 n60 n57 NETTRAN_DUMMY_9538 NETTRAN_DUMMY_9539 AOI21_X1 
XU67 n59 n57 n138 NETTRAN_DUMMY_9540 NETTRAN_DUMMY_9541 XOR2_X1 
XU66 n58 n56 n57 n52 NETTRAN_DUMMY_9542 NETTRAN_DUMMY_9543 OAI21_X1 
XU65 B[22] A[22] n53 NETTRAN_DUMMY_9544 NETTRAN_DUMMY_9545 AND2_X1 
XU64 B[22] A[22] n54 NETTRAN_DUMMY_9546 NETTRAN_DUMMY_9547 NOR2_X1 
XU63 n53 n54 n55 NETTRAN_DUMMY_9548 NETTRAN_DUMMY_9549 NOR2_X1 
XU62 n52 n55 n139 NETTRAN_DUMMY_9550 NETTRAN_DUMMY_9551 XOR2_X1 
XU61 B[23] A[23] n48 NETTRAN_DUMMY_9552 NETTRAN_DUMMY_9553 NOR2_X1 
XU60 B[23] A[23] n50 NETTRAN_DUMMY_9554 NETTRAN_DUMMY_9555 NAND2_X1 
XU59 n8 n50 n51 NETTRAN_DUMMY_9556 NETTRAN_DUMMY_9557 NAND2_X1 
XU58 n53 n9 n52 n49 NETTRAN_DUMMY_9558 NETTRAN_DUMMY_9559 AOI21_X1 
XU57 n51 n49 n140 NETTRAN_DUMMY_9560 NETTRAN_DUMMY_9561 XOR2_X1 
XU56 n50 n48 n49 n44 NETTRAN_DUMMY_9562 NETTRAN_DUMMY_9563 OAI21_X1 
XU55 B[24] A[24] n45 NETTRAN_DUMMY_9564 NETTRAN_DUMMY_9565 AND2_X1 
XU54 B[24] A[24] n46 NETTRAN_DUMMY_9566 NETTRAN_DUMMY_9567 NOR2_X1 
XU53 n45 n46 n47 NETTRAN_DUMMY_9568 NETTRAN_DUMMY_9569 NOR2_X1 
XU52 n44 n47 n127 NETTRAN_DUMMY_9570 NETTRAN_DUMMY_9571 XOR2_X1 
XU51 B[25] A[25] n40 NETTRAN_DUMMY_9572 NETTRAN_DUMMY_9573 NOR2_X1 
XU50 B[25] A[25] n42 NETTRAN_DUMMY_9574 NETTRAN_DUMMY_9575 NAND2_X1 
XU49 n6 n42 n43 NETTRAN_DUMMY_9576 NETTRAN_DUMMY_9577 NAND2_X1 
XU48 n45 n7 n44 n41 NETTRAN_DUMMY_9578 NETTRAN_DUMMY_9579 AOI21_X1 
XU47 n43 n41 n128 NETTRAN_DUMMY_9580 NETTRAN_DUMMY_9581 XOR2_X1 
XU46 n42 n40 n41 n36 NETTRAN_DUMMY_9582 NETTRAN_DUMMY_9583 OAI21_X1 
XU45 B[26] A[26] n37 NETTRAN_DUMMY_9584 NETTRAN_DUMMY_9585 AND2_X1 
XU1 n92 SUM[28] NETTRAN_DUMMY_9586 NETTRAN_DUMMY_9587 BUF_X1 
XU103 n110 SUM[22] NETTRAN_DUMMY_9588 NETTRAN_DUMMY_9589 BUF_X1 
XU104 n123 SUM[18] NETTRAN_DUMMY_9590 NETTRAN_DUMMY_9591 BUF_X1 
XU105 n133 n87 NETTRAN_DUMMY_9592 NETTRAN_DUMMY_9593 INV_X1 
XU106 n87 SUM[30] NETTRAN_DUMMY_9594 NETTRAN_DUMMY_9595 INV_X32 
XU107 n91 n89 NETTRAN_DUMMY_9596 NETTRAN_DUMMY_9597 INV_X1 
XU108 n89 SUM[29] NETTRAN_DUMMY_9598 NETTRAN_DUMMY_9599 INV_X8 
XU109 n132 n91 NETTRAN_DUMMY_9600 NETTRAN_DUMMY_9601 BUF_X32 
XU110 n93 n92 NETTRAN_DUMMY_9602 NETTRAN_DUMMY_9603 CLKBUF_X1 
XU111 n131 n93 NETTRAN_DUMMY_9604 NETTRAN_DUMMY_9605 BUF_X32 
XU112 n96 n94 NETTRAN_DUMMY_9606 NETTRAN_DUMMY_9607 INV_X1 
XU113 n94 SUM[27] NETTRAN_DUMMY_9608 NETTRAN_DUMMY_9609 INV_X32 
XU114 n130 n96 NETTRAN_DUMMY_9610 NETTRAN_DUMMY_9611 BUF_X32 
XU115 n99 n97 NETTRAN_DUMMY_9612 NETTRAN_DUMMY_9613 INV_X1 
XU116 n97 SUM[26] NETTRAN_DUMMY_9614 NETTRAN_DUMMY_9615 INV_X8 
XU117 n129 n99 NETTRAN_DUMMY_9616 NETTRAN_DUMMY_9617 BUF_X32 
XU118 n102 n100 NETTRAN_DUMMY_9618 NETTRAN_DUMMY_9619 INV_X1 
XU119 n100 SUM[25] NETTRAN_DUMMY_9620 NETTRAN_DUMMY_9621 INV_X8 
XU120 n128 n102 NETTRAN_DUMMY_9622 NETTRAN_DUMMY_9623 BUF_X32 
XU121 n105 n103 NETTRAN_DUMMY_9624 NETTRAN_DUMMY_9625 INV_X1 
XU122 n103 SUM[24] NETTRAN_DUMMY_9626 NETTRAN_DUMMY_9627 INV_X8 
XU123 n127 n105 NETTRAN_DUMMY_9628 NETTRAN_DUMMY_9629 BUF_X32 
XU124 n108 n106 NETTRAN_DUMMY_9630 NETTRAN_DUMMY_9631 INV_X1 
XU125 n106 SUM[23] NETTRAN_DUMMY_9632 NETTRAN_DUMMY_9633 INV_X8 
XU126 n140 n108 NETTRAN_DUMMY_9634 NETTRAN_DUMMY_9635 BUF_X32 
XU127 n111 n109 NETTRAN_DUMMY_9636 NETTRAN_DUMMY_9637 INV_X1 
XU128 n109 n110 NETTRAN_DUMMY_9638 NETTRAN_DUMMY_9639 INV_X4 
XU129 n139 n111 NETTRAN_DUMMY_9640 NETTRAN_DUMMY_9641 BUF_X32 
XU130 n114 n112 NETTRAN_DUMMY_9642 NETTRAN_DUMMY_9643 INV_X1 
XU131 n112 SUM[21] NETTRAN_DUMMY_9644 NETTRAN_DUMMY_9645 INV_X8 
XU132 n138 n114 NETTRAN_DUMMY_9646 NETTRAN_DUMMY_9647 BUF_X32 
XU133 n117 n115 NETTRAN_DUMMY_9648 NETTRAN_DUMMY_9649 INV_X1 
XU134 n115 n142 NETTRAN_DUMMY_9650 NETTRAN_DUMMY_9651 INV_X8 
XU135 n137 n117 NETTRAN_DUMMY_9652 NETTRAN_DUMMY_9653 BUF_X32 
XU136 n119 n118 NETTRAN_DUMMY_9654 NETTRAN_DUMMY_9655 CLKBUF_X1 
XU137 n136 n119 NETTRAN_DUMMY_9656 NETTRAN_DUMMY_9657 INV_X1 
XU138 n118 SUM[19] NETTRAN_DUMMY_9658 NETTRAN_DUMMY_9659 INV_X32 
XU139 n122 n121 NETTRAN_DUMMY_9660 NETTRAN_DUMMY_9661 CLKBUF_X1 
XU140 n135 n122 NETTRAN_DUMMY_9662 NETTRAN_DUMMY_9663 INV_X1 
XU141 n121 n123 NETTRAN_DUMMY_9664 NETTRAN_DUMMY_9665 INV_X32 
XU142 n125 n124 NETTRAN_DUMMY_9666 NETTRAN_DUMMY_9667 BUF_X1 
XU143 n134 n125 NETTRAN_DUMMY_9668 NETTRAN_DUMMY_9669 INV_X16 
XU144 n124 SUM[17] NETTRAN_DUMMY_9670 NETTRAN_DUMMY_9671 INV_X32 
XU145 n142 SUM[20] NETTRAN_DUMMY_9672 NETTRAN_DUMMY_9673 BUF_X1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW01_add_0 SUM[37] SUM[36] SUM[35] SUM[34] SUM[33] 
+ SUM[32] SUM[31] SUM[30] SUM[29] SUM[28] SUM[27] SUM[26] SUM[25] SUM[24] SUM[23] 
+ SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] SUM[17] SUM[16] SUM[15] SUM[14] SUM[13] 
+ SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] 
+ SUM[1] SUM[0] CI CO B[37] B[36] B[35] B[34] B[33] B[32] B[31] B[30] B[29] B[28] 
+ B[27] B[26] B[25] B[24] B[23] B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] 
+ B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] 
+ A[37] A[36] A[35] A[34] A[33] A[32] A[31] A[30] A[29] A[28] A[27] A[26] A[25] 
+ A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] A[13] A[12] 
+ A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU1_13 A[13] B[13] carry[13] carry[14] SUM[13] NETTRAN_DUMMY_9674 NETTRAN_DUMMY_9675 FA_X1 
XU1_14 A[14] B[14] carry[14] carry[15] SUM[14] NETTRAN_DUMMY_9676 NETTRAN_DUMMY_9677 FA_X1 
XU1_15 A[15] B[15] carry[15] carry[16] SUM[15] NETTRAN_DUMMY_9678 NETTRAN_DUMMY_9679 FA_X1 
XU1_16 A[16] B[16] carry[16] carry[17] SUM[16] NETTRAN_DUMMY_9680 NETTRAN_DUMMY_9681 FA_X1 
XU1_17 A[17] B[17] carry[17] carry[18] SUM[17] NETTRAN_DUMMY_9682 NETTRAN_DUMMY_9683 FA_X1 
XU1_18 A[18] B[18] carry[18] carry[19] SUM[18] NETTRAN_DUMMY_9684 NETTRAN_DUMMY_9685 FA_X1 
XU1_19 A[19] B[19] carry[19] carry[20] SUM[19] NETTRAN_DUMMY_9686 NETTRAN_DUMMY_9687 FA_X1 
XU1_20 A[20] B[20] carry[20] carry[21] n75 NETTRAN_DUMMY_9688 NETTRAN_DUMMY_9689 FA_X1 
XU1_21 A[21] B[21] carry[21] carry[22] n76 NETTRAN_DUMMY_9690 NETTRAN_DUMMY_9691 FA_X1 
XU1_22 A[22] B[22] carry[22] carry[23] n77 NETTRAN_DUMMY_9692 NETTRAN_DUMMY_9693 FA_X1 
XU1_23 A[23] B[23] carry[23] carry[24] n78 NETTRAN_DUMMY_9694 NETTRAN_DUMMY_9695 FA_X1 
XU1_24 A[24] B[24] carry[24] carry[25] n79 NETTRAN_DUMMY_9696 NETTRAN_DUMMY_9697 FA_X1 
XU1_25 A[25] B[25] carry[25] carry[26] n80 NETTRAN_DUMMY_9698 NETTRAN_DUMMY_9699 FA_X1 
XU1_26 A[26] B[26] carry[26] carry[27] n81 NETTRAN_DUMMY_9700 NETTRAN_DUMMY_9701 FA_X1 
XU1_27 A[27] B[27] carry[27] carry[28] n82 NETTRAN_DUMMY_9702 NETTRAN_DUMMY_9703 FA_X1 
XU1_28 A[28] B[28] carry[28] carry[29] n67 NETTRAN_DUMMY_9704 NETTRAN_DUMMY_9705 FA_X1 
XU1_29 A[29] B[29] carry[29] carry[30] n68 NETTRAN_DUMMY_9706 NETTRAN_DUMMY_9707 FA_X1 
XU1_30 A[30] B[30] carry[30] carry[31] n69 NETTRAN_DUMMY_9708 NETTRAN_DUMMY_9709 FA_X1 
XU1_31 A[31] B[31] carry[31] carry[32] n70 NETTRAN_DUMMY_9710 NETTRAN_DUMMY_9711 FA_X1 
XU1_32 A[32] B[32] carry[32] carry[33] n71 NETTRAN_DUMMY_9712 NETTRAN_DUMMY_9713 FA_X1 
XU1_33 A[33] B[33] carry[33] carry[34] n72 NETTRAN_DUMMY_9714 NETTRAN_DUMMY_9715 FA_X1 
XU1_34 A[34] B[34] carry[34] carry[35] n73 NETTRAN_DUMMY_9716 NETTRAN_DUMMY_9717 FA_X1 
XU1_35 A[35] B[35] carry[35] carry[36] n74 NETTRAN_DUMMY_9718 NETTRAN_DUMMY_9719 FA_X1 
XU1_36 A[36] B[36] carry[36] carry[37] n65 NETTRAN_DUMMY_9720 NETTRAN_DUMMY_9721 FA_X1 
XU1_37 A[37] B[37] carry[37] NETTRAN_DUMMY_9722 n66 NETTRAN_DUMMY_9723 NETTRAN_DUMMY_9724 FA_X1 
XU2 B[0] A[0] SUM[0] NETTRAN_DUMMY_9725 NETTRAN_DUMMY_9726 XOR2_X1 
XU1 B[0] A[0] n1 NETTRAN_DUMMY_9727 NETTRAN_DUMMY_9728 AND2_X1 
XU1_1 A[1] B[1] n1 carry[2] SUM[1] NETTRAN_DUMMY_9729 NETTRAN_DUMMY_9730 FA_X1 
XU1_2 A[2] B[2] carry[2] carry[3] SUM[2] NETTRAN_DUMMY_9731 NETTRAN_DUMMY_9732 FA_X1 
XU1_3 A[3] B[3] carry[3] carry[4] SUM[3] NETTRAN_DUMMY_9733 NETTRAN_DUMMY_9734 FA_X1 
XU1_4 A[4] B[4] carry[4] carry[5] SUM[4] NETTRAN_DUMMY_9735 NETTRAN_DUMMY_9736 FA_X1 
XU1_5 A[5] B[5] carry[5] carry[6] SUM[5] NETTRAN_DUMMY_9737 NETTRAN_DUMMY_9738 FA_X1 
XU1_6 A[6] B[6] carry[6] carry[7] SUM[6] NETTRAN_DUMMY_9739 NETTRAN_DUMMY_9740 FA_X1 
XU1_7 A[7] B[7] carry[7] carry[8] SUM[7] NETTRAN_DUMMY_9741 NETTRAN_DUMMY_9742 FA_X1 
XU1_8 A[8] B[8] carry[8] carry[9] SUM[8] NETTRAN_DUMMY_9743 NETTRAN_DUMMY_9744 FA_X1 
XU1_9 A[9] B[9] carry[9] carry[10] SUM[9] NETTRAN_DUMMY_9745 NETTRAN_DUMMY_9746 FA_X1 
XU1_10 A[10] B[10] carry[10] carry[11] SUM[10] NETTRAN_DUMMY_9747 NETTRAN_DUMMY_9748 FA_X1 
XU1_11 A[11] B[11] carry[11] carry[12] SUM[11] NETTRAN_DUMMY_9749 NETTRAN_DUMMY_9750 FA_X1 
XU1_12 A[12] B[12] carry[12] carry[13] SUM[12] NETTRAN_DUMMY_9751 NETTRAN_DUMMY_9752 FA_X1 
XU3 n3 n2 NETTRAN_DUMMY_9753 NETTRAN_DUMMY_9754 CLKBUF_X1 
XU4 n66 n3 NETTRAN_DUMMY_9755 NETTRAN_DUMMY_9756 INV_X32 
XU5 n2 SUM[37] NETTRAN_DUMMY_9757 NETTRAN_DUMMY_9758 INV_X32 
XU6 n6 n5 NETTRAN_DUMMY_9759 NETTRAN_DUMMY_9760 CLKBUF_X1 
XU7 n65 n6 NETTRAN_DUMMY_9761 NETTRAN_DUMMY_9762 INV_X32 
XU8 n5 SUM[36] NETTRAN_DUMMY_9763 NETTRAN_DUMMY_9764 INV_X32 
XU9 n11 SUM[35] NETTRAN_DUMMY_9765 NETTRAN_DUMMY_9766 BUF_X1 
XU10 n10 n9 NETTRAN_DUMMY_9767 NETTRAN_DUMMY_9768 CLKBUF_X1 
XU11 n74 n10 NETTRAN_DUMMY_9769 NETTRAN_DUMMY_9770 INV_X32 
XU12 n9 n11 NETTRAN_DUMMY_9771 NETTRAN_DUMMY_9772 INV_X32 
XU13 n13 n12 NETTRAN_DUMMY_9773 NETTRAN_DUMMY_9774 CLKBUF_X1 
XU14 n73 n13 NETTRAN_DUMMY_9775 NETTRAN_DUMMY_9776 INV_X32 
XU15 n12 SUM[34] NETTRAN_DUMMY_9777 NETTRAN_DUMMY_9778 INV_X32 
XU16 n18 SUM[33] NETTRAN_DUMMY_9779 NETTRAN_DUMMY_9780 BUF_X1 
XU17 n17 n16 NETTRAN_DUMMY_9781 NETTRAN_DUMMY_9782 CLKBUF_X1 
XU18 n72 n17 NETTRAN_DUMMY_9783 NETTRAN_DUMMY_9784 INV_X32 
XU19 n16 n18 NETTRAN_DUMMY_9785 NETTRAN_DUMMY_9786 INV_X32 
XU20 n22 SUM[32] NETTRAN_DUMMY_9787 NETTRAN_DUMMY_9788 BUF_X1 
XU21 n21 n20 NETTRAN_DUMMY_9789 NETTRAN_DUMMY_9790 CLKBUF_X1 
XU22 n71 n21 NETTRAN_DUMMY_9791 NETTRAN_DUMMY_9792 INV_X32 
XU23 n20 n22 NETTRAN_DUMMY_9793 NETTRAN_DUMMY_9794 INV_X32 
XU24 n26 SUM[31] NETTRAN_DUMMY_9795 NETTRAN_DUMMY_9796 BUF_X1 
XU25 n25 n24 NETTRAN_DUMMY_9797 NETTRAN_DUMMY_9798 CLKBUF_X1 
XU26 n70 n25 NETTRAN_DUMMY_9799 NETTRAN_DUMMY_9800 INV_X32 
XU27 n24 n26 NETTRAN_DUMMY_9801 NETTRAN_DUMMY_9802 INV_X32 
XU28 n28 n27 NETTRAN_DUMMY_9803 NETTRAN_DUMMY_9804 CLKBUF_X1 
XU29 n69 n28 NETTRAN_DUMMY_9805 NETTRAN_DUMMY_9806 INV_X32 
XU30 n27 SUM[30] NETTRAN_DUMMY_9807 NETTRAN_DUMMY_9808 INV_X32 
XU31 n31 n30 NETTRAN_DUMMY_9809 NETTRAN_DUMMY_9810 CLKBUF_X1 
XU32 n68 n31 NETTRAN_DUMMY_9811 NETTRAN_DUMMY_9812 INV_X32 
XU33 n30 SUM[29] NETTRAN_DUMMY_9813 NETTRAN_DUMMY_9814 INV_X32 
XU34 n34 n33 NETTRAN_DUMMY_9815 NETTRAN_DUMMY_9816 CLKBUF_X1 
XU35 n67 n34 NETTRAN_DUMMY_9817 NETTRAN_DUMMY_9818 INV_X32 
XU36 n33 SUM[28] NETTRAN_DUMMY_9819 NETTRAN_DUMMY_9820 INV_X32 
XU37 n37 n36 NETTRAN_DUMMY_9821 NETTRAN_DUMMY_9822 CLKBUF_X1 
XU38 n82 n37 NETTRAN_DUMMY_9823 NETTRAN_DUMMY_9824 INV_X32 
XU39 n36 SUM[27] NETTRAN_DUMMY_9825 NETTRAN_DUMMY_9826 INV_X32 
XU40 n40 n39 NETTRAN_DUMMY_9827 NETTRAN_DUMMY_9828 CLKBUF_X1 
XU41 n81 n40 NETTRAN_DUMMY_9829 NETTRAN_DUMMY_9830 INV_X32 
XU42 n39 SUM[26] NETTRAN_DUMMY_9831 NETTRAN_DUMMY_9832 INV_X32 
XU43 n43 n42 NETTRAN_DUMMY_9833 NETTRAN_DUMMY_9834 CLKBUF_X1 
XU44 n80 n43 NETTRAN_DUMMY_9835 NETTRAN_DUMMY_9836 INV_X32 
XU45 n42 SUM[25] NETTRAN_DUMMY_9837 NETTRAN_DUMMY_9838 INV_X32 
XU46 n48 SUM[24] NETTRAN_DUMMY_9839 NETTRAN_DUMMY_9840 BUF_X1 
XU47 n47 n46 NETTRAN_DUMMY_9841 NETTRAN_DUMMY_9842 CLKBUF_X1 
XU48 n79 n47 NETTRAN_DUMMY_9843 NETTRAN_DUMMY_9844 INV_X32 
XU49 n46 n48 NETTRAN_DUMMY_9845 NETTRAN_DUMMY_9846 INV_X32 
XU50 n52 SUM[23] NETTRAN_DUMMY_9847 NETTRAN_DUMMY_9848 BUF_X1 
XU51 n51 n50 NETTRAN_DUMMY_9849 NETTRAN_DUMMY_9850 CLKBUF_X1 
XU52 n78 n51 NETTRAN_DUMMY_9851 NETTRAN_DUMMY_9852 INV_X32 
XU53 n50 n52 NETTRAN_DUMMY_9853 NETTRAN_DUMMY_9854 INV_X32 
XU54 n56 SUM[22] NETTRAN_DUMMY_9855 NETTRAN_DUMMY_9856 BUF_X1 
XU55 n55 n54 NETTRAN_DUMMY_9857 NETTRAN_DUMMY_9858 CLKBUF_X1 
XU56 n77 n55 NETTRAN_DUMMY_9859 NETTRAN_DUMMY_9860 INV_X32 
XU57 n54 n56 NETTRAN_DUMMY_9861 NETTRAN_DUMMY_9862 INV_X32 
XU58 n60 SUM[21] NETTRAN_DUMMY_9863 NETTRAN_DUMMY_9864 BUF_X1 
XU59 n59 n58 NETTRAN_DUMMY_9865 NETTRAN_DUMMY_9866 CLKBUF_X1 
XU60 n76 n59 NETTRAN_DUMMY_9867 NETTRAN_DUMMY_9868 INV_X32 
XU61 n58 n60 NETTRAN_DUMMY_9869 NETTRAN_DUMMY_9870 INV_X32 
XU62 n64 SUM[20] NETTRAN_DUMMY_9871 NETTRAN_DUMMY_9872 BUF_X1 
XU63 n63 n62 NETTRAN_DUMMY_9873 NETTRAN_DUMMY_9874 CLKBUF_X1 
XU64 n75 n63 NETTRAN_DUMMY_9875 NETTRAN_DUMMY_9876 INV_X32 
XU65 n62 n64 NETTRAN_DUMMY_9877 NETTRAN_DUMMY_9878 INV_X32 
.ENDS

.SUBCKT gng_interp_DW01_inc_0 SUM[15] SUM[14] SUM[13] SUM[12] SUM[11] SUM[10] SUM[9] 
+ SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] A[15] A[14] A[13] 
+ A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU1_1_7 A[7] carry[7] carry[8] SUM[7] NETTRAN_DUMMY_9879 NETTRAN_DUMMY_9880 HA_X1 
XU1_1_6 A[6] carry[6] carry[7] SUM[6] NETTRAN_DUMMY_9881 NETTRAN_DUMMY_9882 HA_X1 
XU1_1_5 A[5] carry[5] carry[6] SUM[5] NETTRAN_DUMMY_9883 NETTRAN_DUMMY_9884 HA_X1 
XU1_1_4 A[4] carry[4] carry[5] SUM[4] NETTRAN_DUMMY_9885 NETTRAN_DUMMY_9886 HA_X1 
XU1_1_3 A[3] carry[3] carry[4] SUM[3] NETTRAN_DUMMY_9887 NETTRAN_DUMMY_9888 HA_X1 
XU1_1_2 A[2] carry[2] carry[3] SUM[2] NETTRAN_DUMMY_9889 NETTRAN_DUMMY_9890 HA_X1 
XU1_1_1 A[1] A[0] carry[2] SUM[1] NETTRAN_DUMMY_9891 NETTRAN_DUMMY_9892 HA_X1 
XU1 carry[15] SUM[15] NETTRAN_DUMMY_9893 NETTRAN_DUMMY_9894 INV_X1 
XU1_1_14 A[14] carry[14] carry[15] SUM[14] NETTRAN_DUMMY_9895 NETTRAN_DUMMY_9896 HA_X1 
XU1_1_13 A[13] carry[13] carry[14] SUM[13] NETTRAN_DUMMY_9897 NETTRAN_DUMMY_9898 HA_X1 
XU1_1_12 A[12] carry[12] carry[13] SUM[12] NETTRAN_DUMMY_9899 NETTRAN_DUMMY_9900 HA_X1 
XU1_1_11 A[11] carry[11] carry[12] SUM[11] NETTRAN_DUMMY_9901 NETTRAN_DUMMY_9902 HA_X1 
XU1_1_10 A[10] carry[10] carry[11] SUM[10] NETTRAN_DUMMY_9903 NETTRAN_DUMMY_9904 HA_X1 
XU1_1_9 A[9] carry[9] carry[10] SUM[9] NETTRAN_DUMMY_9905 NETTRAN_DUMMY_9906 HA_X1 
XU1_1_8 A[8] carry[8] carry[9] SUM[8] NETTRAN_DUMMY_9907 NETTRAN_DUMMY_9908 HA_X1 
.ENDS

.SUBCKT gng_interp_DW01_add_1 SUM[17] SUM[16] SUM[15] SUM[14] SUM[13] SUM[12] SUM[11] 
+ SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
+ CI CO B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] 
+ B[4] B[3] B[2] B[1] B[0] A[17] A[16] A[15] A[14] A[13] A[12] A[11] A[10] A[9] 
+ A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU4 A[0] B[0] A[1] B[1] n3 NETTRAN_DUMMY_9909 NETTRAN_DUMMY_9910 OAI211_X1 
XU3 n3 n2 n1 carry[2] NETTRAN_DUMMY_9911 NETTRAN_DUMMY_9912 OAI21_X1 
XU2 B[1] n1 NETTRAN_DUMMY_9913 NETTRAN_DUMMY_9914 INV_X1 
XU1 A[1] n2 NETTRAN_DUMMY_9915 NETTRAN_DUMMY_9916 INV_X1 
XU1_2 A[2] B[2] carry[2] carry[3] n74 NETTRAN_DUMMY_9917 NETTRAN_DUMMY_9918 FA_X1 
XU1_3 A[3] B[3] carry[3] carry[4] n75 NETTRAN_DUMMY_9919 NETTRAN_DUMMY_9920 FA_X1 
XU1_4 A[4] B[4] carry[4] carry[5] n66 NETTRAN_DUMMY_9921 NETTRAN_DUMMY_9922 FA_X1 
XU1_5 A[5] B[5] carry[5] carry[6] n67 NETTRAN_DUMMY_9923 NETTRAN_DUMMY_9924 FA_X1 
XU1_6 A[6] B[6] carry[6] carry[7] n68 NETTRAN_DUMMY_9925 NETTRAN_DUMMY_9926 FA_X1 
XU1_7 A[7] B[7] carry[7] carry[8] n69 NETTRAN_DUMMY_9927 NETTRAN_DUMMY_9928 FA_X1 
XU1_8 A[8] B[8] carry[8] carry[9] n70 NETTRAN_DUMMY_9929 NETTRAN_DUMMY_9930 FA_X1 
XU1_9 A[9] B[9] carry[9] carry[10] n71 NETTRAN_DUMMY_9931 NETTRAN_DUMMY_9932 FA_X1 
XU1_10 A[10] B[10] carry[10] carry[11] n72 NETTRAN_DUMMY_9933 NETTRAN_DUMMY_9934 FA_X1 
XU1_11 A[11] B[11] carry[11] carry[12] n73 NETTRAN_DUMMY_9935 NETTRAN_DUMMY_9936 FA_X1 
XU1_12 A[12] B[12] carry[12] carry[13] n60 NETTRAN_DUMMY_9937 NETTRAN_DUMMY_9938 FA_X1 
XU1_13 A[13] B[13] carry[13] carry[14] n61 NETTRAN_DUMMY_9939 NETTRAN_DUMMY_9940 FA_X1 
XU1_14 A[14] B[14] carry[14] carry[15] n62 NETTRAN_DUMMY_9941 NETTRAN_DUMMY_9942 FA_X1 
XU1_15 A[15] B[15] carry[15] carry[16] n63 NETTRAN_DUMMY_9943 NETTRAN_DUMMY_9944 FA_X1 
XU1_16 A[16] B[16] carry[16] carry[17] n64 NETTRAN_DUMMY_9945 NETTRAN_DUMMY_9946 FA_X1 
XU1_17 A[17] B[17] carry[17] NETTRAN_DUMMY_9947 n65 NETTRAN_DUMMY_9948 NETTRAN_DUMMY_9949 FA_X1 
XU5 n7 SUM[17] NETTRAN_DUMMY_9950 NETTRAN_DUMMY_9951 BUF_X1 
XU6 n6 n5 NETTRAN_DUMMY_9952 NETTRAN_DUMMY_9953 CLKBUF_X1 
XU7 n65 n6 NETTRAN_DUMMY_9954 NETTRAN_DUMMY_9955 INV_X32 
XU8 n5 n7 NETTRAN_DUMMY_9956 NETTRAN_DUMMY_9957 INV_X32 
XU9 n11 SUM[16] NETTRAN_DUMMY_9958 NETTRAN_DUMMY_9959 BUF_X1 
XU10 n10 n9 NETTRAN_DUMMY_9960 NETTRAN_DUMMY_9961 CLKBUF_X1 
XU11 n64 n10 NETTRAN_DUMMY_9962 NETTRAN_DUMMY_9963 INV_X32 
XU12 n9 n11 NETTRAN_DUMMY_9964 NETTRAN_DUMMY_9965 INV_X32 
XU13 n15 SUM[15] NETTRAN_DUMMY_9966 NETTRAN_DUMMY_9967 BUF_X1 
XU14 n14 n13 NETTRAN_DUMMY_9968 NETTRAN_DUMMY_9969 CLKBUF_X1 
XU15 n63 n14 NETTRAN_DUMMY_9970 NETTRAN_DUMMY_9971 INV_X32 
XU16 n13 n15 NETTRAN_DUMMY_9972 NETTRAN_DUMMY_9973 INV_X32 
XU17 n62 n16 NETTRAN_DUMMY_9974 NETTRAN_DUMMY_9975 CLKBUF_X1 
XU18 n18 n17 NETTRAN_DUMMY_9976 NETTRAN_DUMMY_9977 CLKBUF_X1 
XU19 n16 n18 NETTRAN_DUMMY_9978 NETTRAN_DUMMY_9979 INV_X32 
XU20 n17 SUM[14] NETTRAN_DUMMY_9980 NETTRAN_DUMMY_9981 INV_X32 
XU21 n23 SUM[13] NETTRAN_DUMMY_9982 NETTRAN_DUMMY_9983 CLKBUF_X1 
XU22 n22 n21 NETTRAN_DUMMY_9984 NETTRAN_DUMMY_9985 CLKBUF_X1 
XU23 n61 n22 NETTRAN_DUMMY_9986 NETTRAN_DUMMY_9987 INV_X32 
XU24 n21 n23 NETTRAN_DUMMY_9988 NETTRAN_DUMMY_9989 INV_X32 
XU25 n27 SUM[12] NETTRAN_DUMMY_9990 NETTRAN_DUMMY_9991 BUF_X1 
XU26 n26 n25 NETTRAN_DUMMY_9992 NETTRAN_DUMMY_9993 CLKBUF_X1 
XU27 n60 n26 NETTRAN_DUMMY_9994 NETTRAN_DUMMY_9995 INV_X32 
XU28 n25 n27 NETTRAN_DUMMY_9996 NETTRAN_DUMMY_9997 INV_X32 
XU29 n73 n28 NETTRAN_DUMMY_9998 NETTRAN_DUMMY_9999 CLKBUF_X1 
XU30 n30 n29 NETTRAN_DUMMY_10000 NETTRAN_DUMMY_10001 CLKBUF_X1 
XU31 n28 n30 NETTRAN_DUMMY_10002 NETTRAN_DUMMY_10003 INV_X32 
XU32 n29 SUM[11] NETTRAN_DUMMY_10004 NETTRAN_DUMMY_10005 INV_X32 
XU33 n33 n32 NETTRAN_DUMMY_10006 NETTRAN_DUMMY_10007 CLKBUF_X1 
XU34 n72 n33 NETTRAN_DUMMY_10008 NETTRAN_DUMMY_10009 INV_X32 
XU35 n32 SUM[10] NETTRAN_DUMMY_10010 NETTRAN_DUMMY_10011 INV_X32 
XU36 n36 n35 NETTRAN_DUMMY_10012 NETTRAN_DUMMY_10013 BUF_X1 
XU37 n71 n36 NETTRAN_DUMMY_10014 NETTRAN_DUMMY_10015 INV_X32 
XU38 n35 SUM[9] NETTRAN_DUMMY_10016 NETTRAN_DUMMY_10017 INV_X32 
XU39 n39 n38 NETTRAN_DUMMY_10018 NETTRAN_DUMMY_10019 BUF_X1 
XU40 n70 n39 NETTRAN_DUMMY_10020 NETTRAN_DUMMY_10021 INV_X32 
XU41 n38 SUM[8] NETTRAN_DUMMY_10022 NETTRAN_DUMMY_10023 INV_X32 
XU42 n42 n41 NETTRAN_DUMMY_10024 NETTRAN_DUMMY_10025 CLKBUF_X1 
XU43 n69 n42 NETTRAN_DUMMY_10026 NETTRAN_DUMMY_10027 INV_X32 
XU44 n41 SUM[7] NETTRAN_DUMMY_10028 NETTRAN_DUMMY_10029 INV_X16 
XU45 n47 SUM[6] NETTRAN_DUMMY_10030 NETTRAN_DUMMY_10031 BUF_X1 
XU46 n46 n45 NETTRAN_DUMMY_10032 NETTRAN_DUMMY_10033 CLKBUF_X1 
XU47 n68 n46 NETTRAN_DUMMY_10034 NETTRAN_DUMMY_10035 INV_X32 
XU48 n45 n47 NETTRAN_DUMMY_10036 NETTRAN_DUMMY_10037 INV_X32 
XU49 n49 n48 NETTRAN_DUMMY_10038 NETTRAN_DUMMY_10039 CLKBUF_X1 
XU50 n67 n49 NETTRAN_DUMMY_10040 NETTRAN_DUMMY_10041 INV_X32 
XU51 n48 SUM[5] NETTRAN_DUMMY_10042 NETTRAN_DUMMY_10043 INV_X32 
XU52 n52 n51 NETTRAN_DUMMY_10044 NETTRAN_DUMMY_10045 CLKBUF_X1 
XU53 n66 n52 NETTRAN_DUMMY_10046 NETTRAN_DUMMY_10047 INV_X32 
XU54 n51 SUM[4] NETTRAN_DUMMY_10048 NETTRAN_DUMMY_10049 INV_X32 
XU55 n55 n54 NETTRAN_DUMMY_10050 NETTRAN_DUMMY_10051 BUF_X1 
XU56 n75 n55 NETTRAN_DUMMY_10052 NETTRAN_DUMMY_10053 INV_X32 
XU57 n54 SUM[3] NETTRAN_DUMMY_10054 NETTRAN_DUMMY_10055 INV_X32 
XU58 n58 n57 NETTRAN_DUMMY_10056 NETTRAN_DUMMY_10057 BUF_X1 
XU59 n74 n58 NETTRAN_DUMMY_10058 NETTRAN_DUMMY_10059 INV_X32 
XU60 n57 SUM[2] NETTRAN_DUMMY_10060 NETTRAN_DUMMY_10061 INV_X32 
.ENDS

.SUBCKT gng_smul_16_18_DW02_mult_0 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] 
+ PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] PRODUCT[1] 
+ PRODUCT[0] TC B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] 
+ B[5] B[4] B[3] B[2] B[1] B[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] 
+ A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XS2_14_3 ab_14__3_ CARRYB_13__3_ SUMB_13__4_ CARRYB_14__3_ SUMB_14__3_ NETTRAN_DUMMY_10062 
+ NETTRAN_DUMMY_10063 FA_X1 
XS2_14_2 ab_14__2_ CARRYB_13__2_ SUMB_13__3_ CARRYB_14__2_ SUMB_14__2_ NETTRAN_DUMMY_10064 
+ NETTRAN_DUMMY_10065 FA_X1 
XS2_14_1 ab_14__1_ CARRYB_13__1_ SUMB_13__2_ CARRYB_14__1_ SUMB_14__1_ NETTRAN_DUMMY_10066 
+ NETTRAN_DUMMY_10067 FA_X1 
XS1_14_0 ab_14__0_ CARRYB_13__0_ SUMB_13__1_ CARRYB_14__0_ PRODUCT[14] NETTRAN_DUMMY_10068 
+ NETTRAN_DUMMY_10069 FA_X1 
XS14_17 n1 n85 ab_15__17_ CARRYB_15__17_ SUMB_15__17_ NETTRAN_DUMMY_10070 NETTRAN_DUMMY_10071 FA_X1 
XS5_16 ab_15__16_ CARRYB_14__16_ ab_14__17_ CARRYB_15__16_ SUMB_15__16_ NETTRAN_DUMMY_10072 
+ NETTRAN_DUMMY_10073 FA_X1 
XS4_15 ab_15__15_ CARRYB_14__15_ SUMB_14__16_ CARRYB_15__15_ SUMB_15__15_ NETTRAN_DUMMY_10074 
+ NETTRAN_DUMMY_10075 FA_X1 
XS4_14 ab_15__14_ CARRYB_14__14_ SUMB_14__15_ CARRYB_15__14_ SUMB_15__14_ NETTRAN_DUMMY_10076 
+ NETTRAN_DUMMY_10077 FA_X1 
XS4_13 ab_15__13_ CARRYB_14__13_ SUMB_14__14_ CARRYB_15__13_ SUMB_15__13_ NETTRAN_DUMMY_10078 
+ NETTRAN_DUMMY_10079 FA_X1 
XS4_12 ab_15__12_ CARRYB_14__12_ SUMB_14__13_ CARRYB_15__12_ SUMB_15__12_ NETTRAN_DUMMY_10080 
+ NETTRAN_DUMMY_10081 FA_X1 
XS4_11 ab_15__11_ CARRYB_14__11_ SUMB_14__12_ CARRYB_15__11_ SUMB_15__11_ NETTRAN_DUMMY_10082 
+ NETTRAN_DUMMY_10083 FA_X1 
XS4_10 ab_15__10_ CARRYB_14__10_ SUMB_14__11_ CARRYB_15__10_ SUMB_15__10_ NETTRAN_DUMMY_10084 
+ NETTRAN_DUMMY_10085 FA_X1 
XS4_9 ab_15__9_ CARRYB_14__9_ SUMB_14__10_ CARRYB_15__9_ SUMB_15__9_ NETTRAN_DUMMY_10086 
+ NETTRAN_DUMMY_10087 FA_X1 
XS4_8 ab_15__8_ CARRYB_14__8_ SUMB_14__9_ CARRYB_15__8_ SUMB_15__8_ NETTRAN_DUMMY_10088 
+ NETTRAN_DUMMY_10089 FA_X1 
XS4_7 ab_15__7_ CARRYB_14__7_ SUMB_14__8_ CARRYB_15__7_ SUMB_15__7_ NETTRAN_DUMMY_10090 
+ NETTRAN_DUMMY_10091 FA_X1 
XS4_6 ab_15__6_ CARRYB_14__6_ SUMB_14__7_ CARRYB_15__6_ SUMB_15__6_ NETTRAN_DUMMY_10092 
+ NETTRAN_DUMMY_10093 FA_X1 
XS4_5 ab_15__5_ CARRYB_14__5_ SUMB_14__6_ CARRYB_15__5_ SUMB_15__5_ NETTRAN_DUMMY_10094 
+ NETTRAN_DUMMY_10095 FA_X1 
XS4_4 ab_15__4_ CARRYB_14__4_ SUMB_14__5_ CARRYB_15__4_ SUMB_15__4_ NETTRAN_DUMMY_10096 
+ NETTRAN_DUMMY_10097 FA_X1 
XS4_3 ab_15__3_ CARRYB_14__3_ SUMB_14__4_ CARRYB_15__3_ SUMB_15__3_ NETTRAN_DUMMY_10098 
+ NETTRAN_DUMMY_10099 FA_X1 
XS4_2 ab_15__2_ CARRYB_14__2_ SUMB_14__3_ CARRYB_15__2_ SUMB_15__2_ NETTRAN_DUMMY_10100 
+ NETTRAN_DUMMY_10101 FA_X1 
XS4_1 ab_15__1_ CARRYB_14__1_ SUMB_14__2_ CARRYB_15__1_ SUMB_15__1_ NETTRAN_DUMMY_10102 
+ NETTRAN_DUMMY_10103 FA_X1 
XS4_0 ab_15__0_ CARRYB_14__0_ SUMB_14__1_ CARRYB_15__0_ SUMB_15__0_ NETTRAN_DUMMY_10104 
+ NETTRAN_DUMMY_10105 FA_X1 
XS14_17_0 B[17] CARRYB_15__1_ SUMB_15__2_ A2_16_ A1_15_ NETTRAN_DUMMY_10106 NETTRAN_DUMMY_10107 FA_X1 
XS2_9_11 ab_9__11_ CARRYB_8__11_ SUMB_8__12_ CARRYB_9__11_ SUMB_9__11_ NETTRAN_DUMMY_10108 
+ NETTRAN_DUMMY_10109 FA_X1 
XS2_9_10 ab_9__10_ CARRYB_8__10_ SUMB_8__11_ CARRYB_9__10_ SUMB_9__10_ NETTRAN_DUMMY_10110 
+ NETTRAN_DUMMY_10111 FA_X1 
XS2_9_9 ab_9__9_ CARRYB_8__9_ SUMB_8__10_ CARRYB_9__9_ SUMB_9__9_ NETTRAN_DUMMY_10112 
+ NETTRAN_DUMMY_10113 FA_X1 
XS2_9_8 ab_9__8_ CARRYB_8__8_ SUMB_8__9_ CARRYB_9__8_ SUMB_9__8_ NETTRAN_DUMMY_10114 
+ NETTRAN_DUMMY_10115 FA_X1 
XS2_9_7 ab_9__7_ CARRYB_8__7_ SUMB_8__8_ CARRYB_9__7_ SUMB_9__7_ NETTRAN_DUMMY_10116 
+ NETTRAN_DUMMY_10117 FA_X1 
XS2_9_6 ab_9__6_ CARRYB_8__6_ SUMB_8__7_ CARRYB_9__6_ SUMB_9__6_ NETTRAN_DUMMY_10118 
+ NETTRAN_DUMMY_10119 FA_X1 
XS2_9_5 ab_9__5_ CARRYB_8__5_ SUMB_8__6_ CARRYB_9__5_ SUMB_9__5_ NETTRAN_DUMMY_10120 
+ NETTRAN_DUMMY_10121 FA_X1 
XS2_9_4 ab_9__4_ CARRYB_8__4_ SUMB_8__5_ CARRYB_9__4_ SUMB_9__4_ NETTRAN_DUMMY_10122 
+ NETTRAN_DUMMY_10123 FA_X1 
XS2_9_3 ab_9__3_ CARRYB_8__3_ SUMB_8__4_ CARRYB_9__3_ SUMB_9__3_ NETTRAN_DUMMY_10124 
+ NETTRAN_DUMMY_10125 FA_X1 
XS2_9_2 ab_9__2_ CARRYB_8__2_ SUMB_8__3_ CARRYB_9__2_ SUMB_9__2_ NETTRAN_DUMMY_10126 
+ NETTRAN_DUMMY_10127 FA_X1 
XS2_9_1 ab_9__1_ CARRYB_8__1_ SUMB_8__2_ CARRYB_9__1_ SUMB_9__1_ NETTRAN_DUMMY_10128 
+ NETTRAN_DUMMY_10129 FA_X1 
XS1_9_0 ab_9__0_ CARRYB_8__0_ SUMB_8__1_ CARRYB_9__0_ PRODUCT[9] NETTRAN_DUMMY_10130 
+ NETTRAN_DUMMY_10131 FA_X1 
XS3_10_16 ab_10__16_ CARRYB_9__16_ ab_9__17_ CARRYB_10__16_ SUMB_10__16_ NETTRAN_DUMMY_10132 
+ NETTRAN_DUMMY_10133 FA_X1 
XS2_10_15 ab_10__15_ CARRYB_9__15_ SUMB_9__16_ CARRYB_10__15_ SUMB_10__15_ NETTRAN_DUMMY_10134 
+ NETTRAN_DUMMY_10135 FA_X1 
XS2_10_14 ab_10__14_ CARRYB_9__14_ SUMB_9__15_ CARRYB_10__14_ SUMB_10__14_ NETTRAN_DUMMY_10136 
+ NETTRAN_DUMMY_10137 FA_X1 
XS2_10_13 ab_10__13_ CARRYB_9__13_ SUMB_9__14_ CARRYB_10__13_ SUMB_10__13_ NETTRAN_DUMMY_10138 
+ NETTRAN_DUMMY_10139 FA_X1 
XS2_10_12 ab_10__12_ CARRYB_9__12_ SUMB_9__13_ CARRYB_10__12_ SUMB_10__12_ NETTRAN_DUMMY_10140 
+ NETTRAN_DUMMY_10141 FA_X1 
XS2_10_11 ab_10__11_ CARRYB_9__11_ SUMB_9__12_ CARRYB_10__11_ SUMB_10__11_ NETTRAN_DUMMY_10142 
+ NETTRAN_DUMMY_10143 FA_X1 
XS2_10_10 ab_10__10_ CARRYB_9__10_ SUMB_9__11_ CARRYB_10__10_ SUMB_10__10_ NETTRAN_DUMMY_10144 
+ NETTRAN_DUMMY_10145 FA_X1 
XS2_10_9 ab_10__9_ CARRYB_9__9_ SUMB_9__10_ CARRYB_10__9_ SUMB_10__9_ NETTRAN_DUMMY_10146 
+ NETTRAN_DUMMY_10147 FA_X1 
XS2_10_8 ab_10__8_ CARRYB_9__8_ SUMB_9__9_ CARRYB_10__8_ SUMB_10__8_ NETTRAN_DUMMY_10148 
+ NETTRAN_DUMMY_10149 FA_X1 
XS2_10_7 ab_10__7_ CARRYB_9__7_ SUMB_9__8_ CARRYB_10__7_ SUMB_10__7_ NETTRAN_DUMMY_10150 
+ NETTRAN_DUMMY_10151 FA_X1 
XS2_10_6 ab_10__6_ CARRYB_9__6_ SUMB_9__7_ CARRYB_10__6_ SUMB_10__6_ NETTRAN_DUMMY_10152 
+ NETTRAN_DUMMY_10153 FA_X1 
XS2_10_5 ab_10__5_ CARRYB_9__5_ SUMB_9__6_ CARRYB_10__5_ SUMB_10__5_ NETTRAN_DUMMY_10154 
+ NETTRAN_DUMMY_10155 FA_X1 
XS2_10_4 ab_10__4_ CARRYB_9__4_ SUMB_9__5_ CARRYB_10__4_ SUMB_10__4_ NETTRAN_DUMMY_10156 
+ NETTRAN_DUMMY_10157 FA_X1 
XS2_10_3 ab_10__3_ CARRYB_9__3_ SUMB_9__4_ CARRYB_10__3_ SUMB_10__3_ NETTRAN_DUMMY_10158 
+ NETTRAN_DUMMY_10159 FA_X1 
XS2_10_2 ab_10__2_ CARRYB_9__2_ SUMB_9__3_ CARRYB_10__2_ SUMB_10__2_ NETTRAN_DUMMY_10160 
+ NETTRAN_DUMMY_10161 FA_X1 
XS2_10_1 ab_10__1_ CARRYB_9__1_ SUMB_9__2_ CARRYB_10__1_ SUMB_10__1_ NETTRAN_DUMMY_10162 
+ NETTRAN_DUMMY_10163 FA_X1 
XS1_10_0 ab_10__0_ CARRYB_9__0_ SUMB_9__1_ CARRYB_10__0_ PRODUCT[10] NETTRAN_DUMMY_10164 
+ NETTRAN_DUMMY_10165 FA_X1 
XS3_11_16 ab_11__16_ CARRYB_10__16_ ab_10__17_ CARRYB_11__16_ SUMB_11__16_ NETTRAN_DUMMY_10166 
+ NETTRAN_DUMMY_10167 FA_X1 
XS2_11_15 ab_11__15_ CARRYB_10__15_ SUMB_10__16_ CARRYB_11__15_ SUMB_11__15_ NETTRAN_DUMMY_10168 
+ NETTRAN_DUMMY_10169 FA_X1 
XS2_11_14 ab_11__14_ CARRYB_10__14_ SUMB_10__15_ CARRYB_11__14_ SUMB_11__14_ NETTRAN_DUMMY_10170 
+ NETTRAN_DUMMY_10171 FA_X1 
XS2_11_13 ab_11__13_ CARRYB_10__13_ SUMB_10__14_ CARRYB_11__13_ SUMB_11__13_ NETTRAN_DUMMY_10172 
+ NETTRAN_DUMMY_10173 FA_X1 
XS2_11_12 ab_11__12_ CARRYB_10__12_ SUMB_10__13_ CARRYB_11__12_ SUMB_11__12_ NETTRAN_DUMMY_10174 
+ NETTRAN_DUMMY_10175 FA_X1 
XS2_11_11 ab_11__11_ CARRYB_10__11_ SUMB_10__12_ CARRYB_11__11_ SUMB_11__11_ NETTRAN_DUMMY_10176 
+ NETTRAN_DUMMY_10177 FA_X1 
XS2_11_10 ab_11__10_ CARRYB_10__10_ SUMB_10__11_ CARRYB_11__10_ SUMB_11__10_ NETTRAN_DUMMY_10178 
+ NETTRAN_DUMMY_10179 FA_X1 
XS2_11_9 ab_11__9_ CARRYB_10__9_ SUMB_10__10_ CARRYB_11__9_ SUMB_11__9_ NETTRAN_DUMMY_10180 
+ NETTRAN_DUMMY_10181 FA_X1 
XS2_11_8 ab_11__8_ CARRYB_10__8_ SUMB_10__9_ CARRYB_11__8_ SUMB_11__8_ NETTRAN_DUMMY_10182 
+ NETTRAN_DUMMY_10183 FA_X1 
XS2_11_7 ab_11__7_ CARRYB_10__7_ SUMB_10__8_ CARRYB_11__7_ SUMB_11__7_ NETTRAN_DUMMY_10184 
+ NETTRAN_DUMMY_10185 FA_X1 
XS2_11_6 ab_11__6_ CARRYB_10__6_ SUMB_10__7_ CARRYB_11__6_ SUMB_11__6_ NETTRAN_DUMMY_10186 
+ NETTRAN_DUMMY_10187 FA_X1 
XS2_11_5 ab_11__5_ CARRYB_10__5_ SUMB_10__6_ CARRYB_11__5_ SUMB_11__5_ NETTRAN_DUMMY_10188 
+ NETTRAN_DUMMY_10189 FA_X1 
XS2_11_4 ab_11__4_ CARRYB_10__4_ SUMB_10__5_ CARRYB_11__4_ SUMB_11__4_ NETTRAN_DUMMY_10190 
+ NETTRAN_DUMMY_10191 FA_X1 
XS2_11_3 ab_11__3_ CARRYB_10__3_ SUMB_10__4_ CARRYB_11__3_ SUMB_11__3_ NETTRAN_DUMMY_10192 
+ NETTRAN_DUMMY_10193 FA_X1 
XS2_11_2 ab_11__2_ CARRYB_10__2_ SUMB_10__3_ CARRYB_11__2_ SUMB_11__2_ NETTRAN_DUMMY_10194 
+ NETTRAN_DUMMY_10195 FA_X1 
XS2_11_1 ab_11__1_ CARRYB_10__1_ SUMB_10__2_ CARRYB_11__1_ SUMB_11__1_ NETTRAN_DUMMY_10196 
+ NETTRAN_DUMMY_10197 FA_X1 
XS1_11_0 ab_11__0_ CARRYB_10__0_ SUMB_10__1_ CARRYB_11__0_ PRODUCT[11] NETTRAN_DUMMY_10198 
+ NETTRAN_DUMMY_10199 FA_X1 
XS3_12_16 ab_12__16_ CARRYB_11__16_ ab_11__17_ CARRYB_12__16_ SUMB_12__16_ NETTRAN_DUMMY_10200 
+ NETTRAN_DUMMY_10201 FA_X1 
XS2_12_15 ab_12__15_ CARRYB_11__15_ SUMB_11__16_ CARRYB_12__15_ SUMB_12__15_ NETTRAN_DUMMY_10202 
+ NETTRAN_DUMMY_10203 FA_X1 
XS2_12_14 ab_12__14_ CARRYB_11__14_ SUMB_11__15_ CARRYB_12__14_ SUMB_12__14_ NETTRAN_DUMMY_10204 
+ NETTRAN_DUMMY_10205 FA_X1 
XS2_12_13 ab_12__13_ CARRYB_11__13_ SUMB_11__14_ CARRYB_12__13_ SUMB_12__13_ NETTRAN_DUMMY_10206 
+ NETTRAN_DUMMY_10207 FA_X1 
XS2_12_12 ab_12__12_ CARRYB_11__12_ SUMB_11__13_ CARRYB_12__12_ SUMB_12__12_ NETTRAN_DUMMY_10208 
+ NETTRAN_DUMMY_10209 FA_X1 
XS2_12_11 ab_12__11_ CARRYB_11__11_ SUMB_11__12_ CARRYB_12__11_ SUMB_12__11_ NETTRAN_DUMMY_10210 
+ NETTRAN_DUMMY_10211 FA_X1 
XS2_12_10 ab_12__10_ CARRYB_11__10_ SUMB_11__11_ CARRYB_12__10_ SUMB_12__10_ NETTRAN_DUMMY_10212 
+ NETTRAN_DUMMY_10213 FA_X1 
XS2_12_9 ab_12__9_ CARRYB_11__9_ SUMB_11__10_ CARRYB_12__9_ SUMB_12__9_ NETTRAN_DUMMY_10214 
+ NETTRAN_DUMMY_10215 FA_X1 
XS2_12_8 ab_12__8_ CARRYB_11__8_ SUMB_11__9_ CARRYB_12__8_ SUMB_12__8_ NETTRAN_DUMMY_10216 
+ NETTRAN_DUMMY_10217 FA_X1 
XS2_12_7 ab_12__7_ CARRYB_11__7_ SUMB_11__8_ CARRYB_12__7_ SUMB_12__7_ NETTRAN_DUMMY_10218 
+ NETTRAN_DUMMY_10219 FA_X1 
XS2_12_6 ab_12__6_ CARRYB_11__6_ SUMB_11__7_ CARRYB_12__6_ SUMB_12__6_ NETTRAN_DUMMY_10220 
+ NETTRAN_DUMMY_10221 FA_X1 
XS2_12_5 ab_12__5_ CARRYB_11__5_ SUMB_11__6_ CARRYB_12__5_ SUMB_12__5_ NETTRAN_DUMMY_10222 
+ NETTRAN_DUMMY_10223 FA_X1 
XS2_12_4 ab_12__4_ CARRYB_11__4_ SUMB_11__5_ CARRYB_12__4_ SUMB_12__4_ NETTRAN_DUMMY_10224 
+ NETTRAN_DUMMY_10225 FA_X1 
XS2_12_3 ab_12__3_ CARRYB_11__3_ SUMB_11__4_ CARRYB_12__3_ SUMB_12__3_ NETTRAN_DUMMY_10226 
+ NETTRAN_DUMMY_10227 FA_X1 
XS2_12_2 ab_12__2_ CARRYB_11__2_ SUMB_11__3_ CARRYB_12__2_ SUMB_12__2_ NETTRAN_DUMMY_10228 
+ NETTRAN_DUMMY_10229 FA_X1 
XS2_12_1 ab_12__1_ CARRYB_11__1_ SUMB_11__2_ CARRYB_12__1_ SUMB_12__1_ NETTRAN_DUMMY_10230 
+ NETTRAN_DUMMY_10231 FA_X1 
XS1_12_0 ab_12__0_ CARRYB_11__0_ SUMB_11__1_ CARRYB_12__0_ PRODUCT[12] NETTRAN_DUMMY_10232 
+ NETTRAN_DUMMY_10233 FA_X1 
XS3_13_16 ab_13__16_ CARRYB_12__16_ ab_12__17_ CARRYB_13__16_ SUMB_13__16_ NETTRAN_DUMMY_10234 
+ NETTRAN_DUMMY_10235 FA_X1 
XS2_13_15 ab_13__15_ CARRYB_12__15_ SUMB_12__16_ CARRYB_13__15_ SUMB_13__15_ NETTRAN_DUMMY_10236 
+ NETTRAN_DUMMY_10237 FA_X1 
XS2_13_14 ab_13__14_ CARRYB_12__14_ SUMB_12__15_ CARRYB_13__14_ SUMB_13__14_ NETTRAN_DUMMY_10238 
+ NETTRAN_DUMMY_10239 FA_X1 
XS2_13_13 ab_13__13_ CARRYB_12__13_ SUMB_12__14_ CARRYB_13__13_ SUMB_13__13_ NETTRAN_DUMMY_10240 
+ NETTRAN_DUMMY_10241 FA_X1 
XS2_13_12 ab_13__12_ CARRYB_12__12_ SUMB_12__13_ CARRYB_13__12_ SUMB_13__12_ NETTRAN_DUMMY_10242 
+ NETTRAN_DUMMY_10243 FA_X1 
XS2_13_11 ab_13__11_ CARRYB_12__11_ SUMB_12__12_ CARRYB_13__11_ SUMB_13__11_ NETTRAN_DUMMY_10244 
+ NETTRAN_DUMMY_10245 FA_X1 
XS2_13_10 ab_13__10_ CARRYB_12__10_ SUMB_12__11_ CARRYB_13__10_ SUMB_13__10_ NETTRAN_DUMMY_10246 
+ NETTRAN_DUMMY_10247 FA_X1 
XS2_13_9 ab_13__9_ CARRYB_12__9_ SUMB_12__10_ CARRYB_13__9_ SUMB_13__9_ NETTRAN_DUMMY_10248 
+ NETTRAN_DUMMY_10249 FA_X1 
XS2_13_8 ab_13__8_ CARRYB_12__8_ SUMB_12__9_ CARRYB_13__8_ SUMB_13__8_ NETTRAN_DUMMY_10250 
+ NETTRAN_DUMMY_10251 FA_X1 
XS2_13_7 ab_13__7_ CARRYB_12__7_ SUMB_12__8_ CARRYB_13__7_ SUMB_13__7_ NETTRAN_DUMMY_10252 
+ NETTRAN_DUMMY_10253 FA_X1 
XS2_13_6 ab_13__6_ CARRYB_12__6_ SUMB_12__7_ CARRYB_13__6_ SUMB_13__6_ NETTRAN_DUMMY_10254 
+ NETTRAN_DUMMY_10255 FA_X1 
XS2_13_5 ab_13__5_ CARRYB_12__5_ SUMB_12__6_ CARRYB_13__5_ SUMB_13__5_ NETTRAN_DUMMY_10256 
+ NETTRAN_DUMMY_10257 FA_X1 
XS2_13_4 ab_13__4_ CARRYB_12__4_ SUMB_12__5_ CARRYB_13__4_ SUMB_13__4_ NETTRAN_DUMMY_10258 
+ NETTRAN_DUMMY_10259 FA_X1 
XS2_13_3 ab_13__3_ CARRYB_12__3_ SUMB_12__4_ CARRYB_13__3_ SUMB_13__3_ NETTRAN_DUMMY_10260 
+ NETTRAN_DUMMY_10261 FA_X1 
XS2_13_2 ab_13__2_ CARRYB_12__2_ SUMB_12__3_ CARRYB_13__2_ SUMB_13__2_ NETTRAN_DUMMY_10262 
+ NETTRAN_DUMMY_10263 FA_X1 
XS2_13_1 ab_13__1_ CARRYB_12__1_ SUMB_12__2_ CARRYB_13__1_ SUMB_13__1_ NETTRAN_DUMMY_10264 
+ NETTRAN_DUMMY_10265 FA_X1 
XS1_13_0 ab_13__0_ CARRYB_12__0_ SUMB_12__1_ CARRYB_13__0_ PRODUCT[13] NETTRAN_DUMMY_10266 
+ NETTRAN_DUMMY_10267 FA_X1 
XS3_14_16 ab_14__16_ CARRYB_13__16_ ab_13__17_ CARRYB_14__16_ SUMB_14__16_ NETTRAN_DUMMY_10268 
+ NETTRAN_DUMMY_10269 FA_X1 
XS2_14_15 ab_14__15_ CARRYB_13__15_ SUMB_13__16_ CARRYB_14__15_ SUMB_14__15_ NETTRAN_DUMMY_10270 
+ NETTRAN_DUMMY_10271 FA_X1 
XS2_14_14 ab_14__14_ CARRYB_13__14_ SUMB_13__15_ CARRYB_14__14_ SUMB_14__14_ NETTRAN_DUMMY_10272 
+ NETTRAN_DUMMY_10273 FA_X1 
XS2_14_13 ab_14__13_ CARRYB_13__13_ SUMB_13__14_ CARRYB_14__13_ SUMB_14__13_ NETTRAN_DUMMY_10274 
+ NETTRAN_DUMMY_10275 FA_X1 
XS2_14_12 ab_14__12_ CARRYB_13__12_ SUMB_13__13_ CARRYB_14__12_ SUMB_14__12_ NETTRAN_DUMMY_10276 
+ NETTRAN_DUMMY_10277 FA_X1 
XS2_14_11 ab_14__11_ CARRYB_13__11_ SUMB_13__12_ CARRYB_14__11_ SUMB_14__11_ NETTRAN_DUMMY_10278 
+ NETTRAN_DUMMY_10279 FA_X1 
XS2_14_10 ab_14__10_ CARRYB_13__10_ SUMB_13__11_ CARRYB_14__10_ SUMB_14__10_ NETTRAN_DUMMY_10280 
+ NETTRAN_DUMMY_10281 FA_X1 
XS2_14_9 ab_14__9_ CARRYB_13__9_ SUMB_13__10_ CARRYB_14__9_ SUMB_14__9_ NETTRAN_DUMMY_10282 
+ NETTRAN_DUMMY_10283 FA_X1 
XS2_14_8 ab_14__8_ CARRYB_13__8_ SUMB_13__9_ CARRYB_14__8_ SUMB_14__8_ NETTRAN_DUMMY_10284 
+ NETTRAN_DUMMY_10285 FA_X1 
XS2_14_7 ab_14__7_ CARRYB_13__7_ SUMB_13__8_ CARRYB_14__7_ SUMB_14__7_ NETTRAN_DUMMY_10286 
+ NETTRAN_DUMMY_10287 FA_X1 
XS2_14_6 ab_14__6_ CARRYB_13__6_ SUMB_13__7_ CARRYB_14__6_ SUMB_14__6_ NETTRAN_DUMMY_10288 
+ NETTRAN_DUMMY_10289 FA_X1 
XS2_14_5 ab_14__5_ CARRYB_13__5_ SUMB_13__6_ CARRYB_14__5_ SUMB_14__5_ NETTRAN_DUMMY_10290 
+ NETTRAN_DUMMY_10291 FA_X1 
XS2_14_4 ab_14__4_ CARRYB_13__4_ SUMB_13__5_ CARRYB_14__4_ SUMB_14__4_ NETTRAN_DUMMY_10292 
+ NETTRAN_DUMMY_10293 FA_X1 
XS2_3_2 ab_3__2_ CARRYB_2__2_ SUMB_2__3_ CARRYB_3__2_ SUMB_3__2_ NETTRAN_DUMMY_10294 
+ NETTRAN_DUMMY_10295 FA_X1 
XS2_3_1 ab_3__1_ CARRYB_2__1_ SUMB_2__2_ CARRYB_3__1_ SUMB_3__1_ NETTRAN_DUMMY_10296 
+ NETTRAN_DUMMY_10297 FA_X1 
XS1_3_0 ab_3__0_ CARRYB_2__0_ SUMB_2__1_ CARRYB_3__0_ PRODUCT[3] NETTRAN_DUMMY_10298 
+ NETTRAN_DUMMY_10299 FA_X1 
XS3_4_16 ab_4__16_ CARRYB_3__16_ ab_3__17_ CARRYB_4__16_ SUMB_4__16_ NETTRAN_DUMMY_10300 
+ NETTRAN_DUMMY_10301 FA_X1 
XS2_4_15 ab_4__15_ CARRYB_3__15_ SUMB_3__16_ CARRYB_4__15_ SUMB_4__15_ NETTRAN_DUMMY_10302 
+ NETTRAN_DUMMY_10303 FA_X1 
XS2_4_14 ab_4__14_ CARRYB_3__14_ SUMB_3__15_ CARRYB_4__14_ SUMB_4__14_ NETTRAN_DUMMY_10304 
+ NETTRAN_DUMMY_10305 FA_X1 
XS2_4_13 ab_4__13_ CARRYB_3__13_ SUMB_3__14_ CARRYB_4__13_ SUMB_4__13_ NETTRAN_DUMMY_10306 
+ NETTRAN_DUMMY_10307 FA_X1 
XS2_4_12 ab_4__12_ CARRYB_3__12_ SUMB_3__13_ CARRYB_4__12_ SUMB_4__12_ NETTRAN_DUMMY_10308 
+ NETTRAN_DUMMY_10309 FA_X1 
XS2_4_11 ab_4__11_ CARRYB_3__11_ SUMB_3__12_ CARRYB_4__11_ SUMB_4__11_ NETTRAN_DUMMY_10310 
+ NETTRAN_DUMMY_10311 FA_X1 
XS2_4_10 ab_4__10_ CARRYB_3__10_ SUMB_3__11_ CARRYB_4__10_ SUMB_4__10_ NETTRAN_DUMMY_10312 
+ NETTRAN_DUMMY_10313 FA_X1 
XS2_4_9 ab_4__9_ CARRYB_3__9_ SUMB_3__10_ CARRYB_4__9_ SUMB_4__9_ NETTRAN_DUMMY_10314 
+ NETTRAN_DUMMY_10315 FA_X1 
XS2_4_8 ab_4__8_ CARRYB_3__8_ SUMB_3__9_ CARRYB_4__8_ SUMB_4__8_ NETTRAN_DUMMY_10316 
+ NETTRAN_DUMMY_10317 FA_X1 
XS2_4_7 ab_4__7_ CARRYB_3__7_ SUMB_3__8_ CARRYB_4__7_ SUMB_4__7_ NETTRAN_DUMMY_10318 
+ NETTRAN_DUMMY_10319 FA_X1 
XS2_4_6 ab_4__6_ CARRYB_3__6_ SUMB_3__7_ CARRYB_4__6_ SUMB_4__6_ NETTRAN_DUMMY_10320 
+ NETTRAN_DUMMY_10321 FA_X1 
XS2_4_5 ab_4__5_ CARRYB_3__5_ SUMB_3__6_ CARRYB_4__5_ SUMB_4__5_ NETTRAN_DUMMY_10322 
+ NETTRAN_DUMMY_10323 FA_X1 
XS2_4_4 ab_4__4_ CARRYB_3__4_ SUMB_3__5_ CARRYB_4__4_ SUMB_4__4_ NETTRAN_DUMMY_10324 
+ NETTRAN_DUMMY_10325 FA_X1 
XS2_4_3 ab_4__3_ CARRYB_3__3_ SUMB_3__4_ CARRYB_4__3_ SUMB_4__3_ NETTRAN_DUMMY_10326 
+ NETTRAN_DUMMY_10327 FA_X1 
XS2_4_2 ab_4__2_ CARRYB_3__2_ SUMB_3__3_ CARRYB_4__2_ SUMB_4__2_ NETTRAN_DUMMY_10328 
+ NETTRAN_DUMMY_10329 FA_X1 
XS2_4_1 ab_4__1_ CARRYB_3__1_ SUMB_3__2_ CARRYB_4__1_ SUMB_4__1_ NETTRAN_DUMMY_10330 
+ NETTRAN_DUMMY_10331 FA_X1 
XS1_4_0 ab_4__0_ CARRYB_3__0_ SUMB_3__1_ CARRYB_4__0_ PRODUCT[4] NETTRAN_DUMMY_10332 
+ NETTRAN_DUMMY_10333 FA_X1 
XS3_5_16 ab_5__16_ CARRYB_4__16_ ab_4__17_ CARRYB_5__16_ SUMB_5__16_ NETTRAN_DUMMY_10334 
+ NETTRAN_DUMMY_10335 FA_X1 
XS2_5_15 ab_5__15_ CARRYB_4__15_ SUMB_4__16_ CARRYB_5__15_ SUMB_5__15_ NETTRAN_DUMMY_10336 
+ NETTRAN_DUMMY_10337 FA_X1 
XS2_5_14 ab_5__14_ CARRYB_4__14_ SUMB_4__15_ CARRYB_5__14_ SUMB_5__14_ NETTRAN_DUMMY_10338 
+ NETTRAN_DUMMY_10339 FA_X1 
XS2_5_13 ab_5__13_ CARRYB_4__13_ SUMB_4__14_ CARRYB_5__13_ SUMB_5__13_ NETTRAN_DUMMY_10340 
+ NETTRAN_DUMMY_10341 FA_X1 
XS2_5_12 ab_5__12_ CARRYB_4__12_ SUMB_4__13_ CARRYB_5__12_ SUMB_5__12_ NETTRAN_DUMMY_10342 
+ NETTRAN_DUMMY_10343 FA_X1 
XS2_5_11 ab_5__11_ CARRYB_4__11_ SUMB_4__12_ CARRYB_5__11_ SUMB_5__11_ NETTRAN_DUMMY_10344 
+ NETTRAN_DUMMY_10345 FA_X1 
XS2_5_10 ab_5__10_ CARRYB_4__10_ SUMB_4__11_ CARRYB_5__10_ SUMB_5__10_ NETTRAN_DUMMY_10346 
+ NETTRAN_DUMMY_10347 FA_X1 
XS2_5_9 ab_5__9_ CARRYB_4__9_ SUMB_4__10_ CARRYB_5__9_ SUMB_5__9_ NETTRAN_DUMMY_10348 
+ NETTRAN_DUMMY_10349 FA_X1 
XS2_5_8 ab_5__8_ CARRYB_4__8_ SUMB_4__9_ CARRYB_5__8_ SUMB_5__8_ NETTRAN_DUMMY_10350 
+ NETTRAN_DUMMY_10351 FA_X1 
XS2_5_7 ab_5__7_ CARRYB_4__7_ SUMB_4__8_ CARRYB_5__7_ SUMB_5__7_ NETTRAN_DUMMY_10352 
+ NETTRAN_DUMMY_10353 FA_X1 
XS2_5_6 ab_5__6_ CARRYB_4__6_ SUMB_4__7_ CARRYB_5__6_ SUMB_5__6_ NETTRAN_DUMMY_10354 
+ NETTRAN_DUMMY_10355 FA_X1 
XS2_5_5 ab_5__5_ CARRYB_4__5_ SUMB_4__6_ CARRYB_5__5_ SUMB_5__5_ NETTRAN_DUMMY_10356 
+ NETTRAN_DUMMY_10357 FA_X1 
XS2_5_4 ab_5__4_ CARRYB_4__4_ SUMB_4__5_ CARRYB_5__4_ SUMB_5__4_ NETTRAN_DUMMY_10358 
+ NETTRAN_DUMMY_10359 FA_X1 
XS2_5_3 ab_5__3_ CARRYB_4__3_ SUMB_4__4_ CARRYB_5__3_ SUMB_5__3_ NETTRAN_DUMMY_10360 
+ NETTRAN_DUMMY_10361 FA_X1 
XS2_5_2 ab_5__2_ CARRYB_4__2_ SUMB_4__3_ CARRYB_5__2_ SUMB_5__2_ NETTRAN_DUMMY_10362 
+ NETTRAN_DUMMY_10363 FA_X1 
XS2_5_1 ab_5__1_ CARRYB_4__1_ SUMB_4__2_ CARRYB_5__1_ SUMB_5__1_ NETTRAN_DUMMY_10364 
+ NETTRAN_DUMMY_10365 FA_X1 
XS1_5_0 ab_5__0_ CARRYB_4__0_ SUMB_4__1_ CARRYB_5__0_ PRODUCT[5] NETTRAN_DUMMY_10366 
+ NETTRAN_DUMMY_10367 FA_X1 
XS3_6_16 ab_6__16_ CARRYB_5__16_ ab_5__17_ CARRYB_6__16_ SUMB_6__16_ NETTRAN_DUMMY_10368 
+ NETTRAN_DUMMY_10369 FA_X1 
XS2_6_15 ab_6__15_ CARRYB_5__15_ SUMB_5__16_ CARRYB_6__15_ SUMB_6__15_ NETTRAN_DUMMY_10370 
+ NETTRAN_DUMMY_10371 FA_X1 
XS2_6_14 ab_6__14_ CARRYB_5__14_ SUMB_5__15_ CARRYB_6__14_ SUMB_6__14_ NETTRAN_DUMMY_10372 
+ NETTRAN_DUMMY_10373 FA_X1 
XS2_6_13 ab_6__13_ CARRYB_5__13_ SUMB_5__14_ CARRYB_6__13_ SUMB_6__13_ NETTRAN_DUMMY_10374 
+ NETTRAN_DUMMY_10375 FA_X1 
XS2_6_12 ab_6__12_ CARRYB_5__12_ SUMB_5__13_ CARRYB_6__12_ SUMB_6__12_ NETTRAN_DUMMY_10376 
+ NETTRAN_DUMMY_10377 FA_X1 
XS2_6_11 ab_6__11_ CARRYB_5__11_ SUMB_5__12_ CARRYB_6__11_ SUMB_6__11_ NETTRAN_DUMMY_10378 
+ NETTRAN_DUMMY_10379 FA_X1 
XS2_6_10 ab_6__10_ CARRYB_5__10_ SUMB_5__11_ CARRYB_6__10_ SUMB_6__10_ NETTRAN_DUMMY_10380 
+ NETTRAN_DUMMY_10381 FA_X1 
XS2_6_9 ab_6__9_ CARRYB_5__9_ SUMB_5__10_ CARRYB_6__9_ SUMB_6__9_ NETTRAN_DUMMY_10382 
+ NETTRAN_DUMMY_10383 FA_X1 
XS2_6_8 ab_6__8_ CARRYB_5__8_ SUMB_5__9_ CARRYB_6__8_ SUMB_6__8_ NETTRAN_DUMMY_10384 
+ NETTRAN_DUMMY_10385 FA_X1 
XS2_6_7 ab_6__7_ CARRYB_5__7_ SUMB_5__8_ CARRYB_6__7_ SUMB_6__7_ NETTRAN_DUMMY_10386 
+ NETTRAN_DUMMY_10387 FA_X1 
XS2_6_6 ab_6__6_ CARRYB_5__6_ SUMB_5__7_ CARRYB_6__6_ SUMB_6__6_ NETTRAN_DUMMY_10388 
+ NETTRAN_DUMMY_10389 FA_X1 
XS2_6_5 ab_6__5_ CARRYB_5__5_ SUMB_5__6_ CARRYB_6__5_ SUMB_6__5_ NETTRAN_DUMMY_10390 
+ NETTRAN_DUMMY_10391 FA_X1 
XS2_6_4 ab_6__4_ CARRYB_5__4_ SUMB_5__5_ CARRYB_6__4_ SUMB_6__4_ NETTRAN_DUMMY_10392 
+ NETTRAN_DUMMY_10393 FA_X1 
XS2_6_3 ab_6__3_ CARRYB_5__3_ SUMB_5__4_ CARRYB_6__3_ SUMB_6__3_ NETTRAN_DUMMY_10394 
+ NETTRAN_DUMMY_10395 FA_X1 
XS2_6_2 ab_6__2_ CARRYB_5__2_ SUMB_5__3_ CARRYB_6__2_ SUMB_6__2_ NETTRAN_DUMMY_10396 
+ NETTRAN_DUMMY_10397 FA_X1 
XS2_6_1 ab_6__1_ CARRYB_5__1_ SUMB_5__2_ CARRYB_6__1_ SUMB_6__1_ NETTRAN_DUMMY_10398 
+ NETTRAN_DUMMY_10399 FA_X1 
XS1_6_0 ab_6__0_ CARRYB_5__0_ SUMB_5__1_ CARRYB_6__0_ PRODUCT[6] NETTRAN_DUMMY_10400 
+ NETTRAN_DUMMY_10401 FA_X1 
XS3_7_16 ab_7__16_ CARRYB_6__16_ ab_6__17_ CARRYB_7__16_ SUMB_7__16_ NETTRAN_DUMMY_10402 
+ NETTRAN_DUMMY_10403 FA_X1 
XS2_7_15 ab_7__15_ CARRYB_6__15_ SUMB_6__16_ CARRYB_7__15_ SUMB_7__15_ NETTRAN_DUMMY_10404 
+ NETTRAN_DUMMY_10405 FA_X1 
XS2_7_14 ab_7__14_ CARRYB_6__14_ SUMB_6__15_ CARRYB_7__14_ SUMB_7__14_ NETTRAN_DUMMY_10406 
+ NETTRAN_DUMMY_10407 FA_X1 
XS2_7_13 ab_7__13_ CARRYB_6__13_ SUMB_6__14_ CARRYB_7__13_ SUMB_7__13_ NETTRAN_DUMMY_10408 
+ NETTRAN_DUMMY_10409 FA_X1 
XS2_7_12 ab_7__12_ CARRYB_6__12_ SUMB_6__13_ CARRYB_7__12_ SUMB_7__12_ NETTRAN_DUMMY_10410 
+ NETTRAN_DUMMY_10411 FA_X1 
XS2_7_11 ab_7__11_ CARRYB_6__11_ SUMB_6__12_ CARRYB_7__11_ SUMB_7__11_ NETTRAN_DUMMY_10412 
+ NETTRAN_DUMMY_10413 FA_X1 
XS2_7_10 ab_7__10_ CARRYB_6__10_ SUMB_6__11_ CARRYB_7__10_ SUMB_7__10_ NETTRAN_DUMMY_10414 
+ NETTRAN_DUMMY_10415 FA_X1 
XS2_7_9 ab_7__9_ CARRYB_6__9_ SUMB_6__10_ CARRYB_7__9_ SUMB_7__9_ NETTRAN_DUMMY_10416 
+ NETTRAN_DUMMY_10417 FA_X1 
XS2_7_8 ab_7__8_ CARRYB_6__8_ SUMB_6__9_ CARRYB_7__8_ SUMB_7__8_ NETTRAN_DUMMY_10418 
+ NETTRAN_DUMMY_10419 FA_X1 
XS2_7_7 ab_7__7_ CARRYB_6__7_ SUMB_6__8_ CARRYB_7__7_ SUMB_7__7_ NETTRAN_DUMMY_10420 
+ NETTRAN_DUMMY_10421 FA_X1 
XS2_7_6 ab_7__6_ CARRYB_6__6_ SUMB_6__7_ CARRYB_7__6_ SUMB_7__6_ NETTRAN_DUMMY_10422 
+ NETTRAN_DUMMY_10423 FA_X1 
XS2_7_5 ab_7__5_ CARRYB_6__5_ SUMB_6__6_ CARRYB_7__5_ SUMB_7__5_ NETTRAN_DUMMY_10424 
+ NETTRAN_DUMMY_10425 FA_X1 
XS2_7_4 ab_7__4_ CARRYB_6__4_ SUMB_6__5_ CARRYB_7__4_ SUMB_7__4_ NETTRAN_DUMMY_10426 
+ NETTRAN_DUMMY_10427 FA_X1 
XS2_7_3 ab_7__3_ CARRYB_6__3_ SUMB_6__4_ CARRYB_7__3_ SUMB_7__3_ NETTRAN_DUMMY_10428 
+ NETTRAN_DUMMY_10429 FA_X1 
XS2_7_2 ab_7__2_ CARRYB_6__2_ SUMB_6__3_ CARRYB_7__2_ SUMB_7__2_ NETTRAN_DUMMY_10430 
+ NETTRAN_DUMMY_10431 FA_X1 
XS2_7_1 ab_7__1_ CARRYB_6__1_ SUMB_6__2_ CARRYB_7__1_ SUMB_7__1_ NETTRAN_DUMMY_10432 
+ NETTRAN_DUMMY_10433 FA_X1 
XS1_7_0 ab_7__0_ CARRYB_6__0_ SUMB_6__1_ CARRYB_7__0_ PRODUCT[7] NETTRAN_DUMMY_10434 
+ NETTRAN_DUMMY_10435 FA_X1 
XS3_8_16 ab_8__16_ CARRYB_7__16_ ab_7__17_ CARRYB_8__16_ SUMB_8__16_ NETTRAN_DUMMY_10436 
+ NETTRAN_DUMMY_10437 FA_X1 
XS2_8_15 ab_8__15_ CARRYB_7__15_ SUMB_7__16_ CARRYB_8__15_ SUMB_8__15_ NETTRAN_DUMMY_10438 
+ NETTRAN_DUMMY_10439 FA_X1 
XS2_8_14 ab_8__14_ CARRYB_7__14_ SUMB_7__15_ CARRYB_8__14_ SUMB_8__14_ NETTRAN_DUMMY_10440 
+ NETTRAN_DUMMY_10441 FA_X1 
XS2_8_13 ab_8__13_ CARRYB_7__13_ SUMB_7__14_ CARRYB_8__13_ SUMB_8__13_ NETTRAN_DUMMY_10442 
+ NETTRAN_DUMMY_10443 FA_X1 
XS2_8_12 ab_8__12_ CARRYB_7__12_ SUMB_7__13_ CARRYB_8__12_ SUMB_8__12_ NETTRAN_DUMMY_10444 
+ NETTRAN_DUMMY_10445 FA_X1 
XS2_8_11 ab_8__11_ CARRYB_7__11_ SUMB_7__12_ CARRYB_8__11_ SUMB_8__11_ NETTRAN_DUMMY_10446 
+ NETTRAN_DUMMY_10447 FA_X1 
XS2_8_10 ab_8__10_ CARRYB_7__10_ SUMB_7__11_ CARRYB_8__10_ SUMB_8__10_ NETTRAN_DUMMY_10448 
+ NETTRAN_DUMMY_10449 FA_X1 
XS2_8_9 ab_8__9_ CARRYB_7__9_ SUMB_7__10_ CARRYB_8__9_ SUMB_8__9_ NETTRAN_DUMMY_10450 
+ NETTRAN_DUMMY_10451 FA_X1 
XS2_8_8 ab_8__8_ CARRYB_7__8_ SUMB_7__9_ CARRYB_8__8_ SUMB_8__8_ NETTRAN_DUMMY_10452 
+ NETTRAN_DUMMY_10453 FA_X1 
XS2_8_7 ab_8__7_ CARRYB_7__7_ SUMB_7__8_ CARRYB_8__7_ SUMB_8__7_ NETTRAN_DUMMY_10454 
+ NETTRAN_DUMMY_10455 FA_X1 
XS2_8_6 ab_8__6_ CARRYB_7__6_ SUMB_7__7_ CARRYB_8__6_ SUMB_8__6_ NETTRAN_DUMMY_10456 
+ NETTRAN_DUMMY_10457 FA_X1 
XS2_8_5 ab_8__5_ CARRYB_7__5_ SUMB_7__6_ CARRYB_8__5_ SUMB_8__5_ NETTRAN_DUMMY_10458 
+ NETTRAN_DUMMY_10459 FA_X1 
XS2_8_4 ab_8__4_ CARRYB_7__4_ SUMB_7__5_ CARRYB_8__4_ SUMB_8__4_ NETTRAN_DUMMY_10460 
+ NETTRAN_DUMMY_10461 FA_X1 
XS2_8_3 ab_8__3_ CARRYB_7__3_ SUMB_7__4_ CARRYB_8__3_ SUMB_8__3_ NETTRAN_DUMMY_10462 
+ NETTRAN_DUMMY_10463 FA_X1 
XS2_8_2 ab_8__2_ CARRYB_7__2_ SUMB_7__3_ CARRYB_8__2_ SUMB_8__2_ NETTRAN_DUMMY_10464 
+ NETTRAN_DUMMY_10465 FA_X1 
XS2_8_1 ab_8__1_ CARRYB_7__1_ SUMB_7__2_ CARRYB_8__1_ SUMB_8__1_ NETTRAN_DUMMY_10466 
+ NETTRAN_DUMMY_10467 FA_X1 
XS1_8_0 ab_8__0_ CARRYB_7__0_ SUMB_7__1_ CARRYB_8__0_ PRODUCT[8] NETTRAN_DUMMY_10468 
+ NETTRAN_DUMMY_10469 FA_X1 
XS3_9_16 ab_9__16_ CARRYB_8__16_ ab_8__17_ CARRYB_9__16_ SUMB_9__16_ NETTRAN_DUMMY_10470 
+ NETTRAN_DUMMY_10471 FA_X1 
XS2_9_15 ab_9__15_ CARRYB_8__15_ SUMB_8__16_ CARRYB_9__15_ SUMB_9__15_ NETTRAN_DUMMY_10472 
+ NETTRAN_DUMMY_10473 FA_X1 
XS2_9_14 ab_9__14_ CARRYB_8__14_ SUMB_8__15_ CARRYB_9__14_ SUMB_9__14_ NETTRAN_DUMMY_10474 
+ NETTRAN_DUMMY_10475 FA_X1 
XS2_9_13 ab_9__13_ CARRYB_8__13_ SUMB_8__14_ CARRYB_9__13_ SUMB_9__13_ NETTRAN_DUMMY_10476 
+ NETTRAN_DUMMY_10477 FA_X1 
XS2_9_12 ab_9__12_ CARRYB_8__12_ SUMB_8__13_ CARRYB_9__12_ SUMB_9__12_ NETTRAN_DUMMY_10478 
+ NETTRAN_DUMMY_10479 FA_X1 
XU63 CARRYB_15__5_ SUMB_15__6_ n62 NETTRAN_DUMMY_10480 NETTRAN_DUMMY_10481 XOR2_X1 
XU62 CARRYB_15__15_ SUMB_15__16_ n61 NETTRAN_DUMMY_10482 NETTRAN_DUMMY_10483 AND2_X1 
XU61 CARRYB_15__14_ SUMB_15__15_ n60 NETTRAN_DUMMY_10484 NETTRAN_DUMMY_10485 AND2_X1 
XU60 CARRYB_15__13_ SUMB_15__14_ n59 NETTRAN_DUMMY_10486 NETTRAN_DUMMY_10487 AND2_X1 
XU59 CARRYB_15__12_ SUMB_15__13_ n58 NETTRAN_DUMMY_10488 NETTRAN_DUMMY_10489 AND2_X1 
XU58 CARRYB_15__11_ SUMB_15__12_ n57 NETTRAN_DUMMY_10490 NETTRAN_DUMMY_10491 AND2_X1 
XU57 CARRYB_15__10_ SUMB_15__11_ n56 NETTRAN_DUMMY_10492 NETTRAN_DUMMY_10493 AND2_X1 
XU56 CARRYB_15__9_ SUMB_15__10_ n55 NETTRAN_DUMMY_10494 NETTRAN_DUMMY_10495 AND2_X1 
XU55 CARRYB_15__8_ SUMB_15__9_ n54 NETTRAN_DUMMY_10496 NETTRAN_DUMMY_10497 AND2_X1 
XU54 CARRYB_15__7_ SUMB_15__8_ n53 NETTRAN_DUMMY_10498 NETTRAN_DUMMY_10499 AND2_X1 
XU53 CARRYB_15__6_ SUMB_15__7_ n52 NETTRAN_DUMMY_10500 NETTRAN_DUMMY_10501 AND2_X1 
XU52 CARRYB_15__5_ SUMB_15__6_ n51 NETTRAN_DUMMY_10502 NETTRAN_DUMMY_10503 AND2_X1 
XU51 CARRYB_15__4_ SUMB_15__5_ n50 NETTRAN_DUMMY_10504 NETTRAN_DUMMY_10505 AND2_X1 
XU50 CARRYB_15__16_ SUMB_15__17_ n49 NETTRAN_DUMMY_10506 NETTRAN_DUMMY_10507 AND2_X1 
XU49 CARRYB_15__16_ SUMB_15__17_ n48 NETTRAN_DUMMY_10508 NETTRAN_DUMMY_10509 XOR2_X1 
XU48 CARRYB_15__14_ SUMB_15__15_ n47 NETTRAN_DUMMY_10510 NETTRAN_DUMMY_10511 XOR2_X1 
XU47 CARRYB_15__12_ SUMB_15__13_ n46 NETTRAN_DUMMY_10512 NETTRAN_DUMMY_10513 XOR2_X1 
XU46 CARRYB_15__10_ SUMB_15__11_ n45 NETTRAN_DUMMY_10514 NETTRAN_DUMMY_10515 XOR2_X1 
XU45 CARRYB_15__8_ SUMB_15__9_ n44 NETTRAN_DUMMY_10516 NETTRAN_DUMMY_10517 XOR2_X1 
XU44 CARRYB_15__6_ SUMB_15__7_ n43 NETTRAN_DUMMY_10518 NETTRAN_DUMMY_10519 XOR2_X1 
XU43 CARRYB_15__3_ SUMB_15__4_ n42 NETTRAN_DUMMY_10520 NETTRAN_DUMMY_10521 XOR2_X1 
XU42 CARRYB_15__3_ SUMB_15__4_ n41 NETTRAN_DUMMY_10522 NETTRAN_DUMMY_10523 AND2_X1 
XU41 CARRYB_15__2_ SUMB_15__3_ n40 NETTRAN_DUMMY_10524 NETTRAN_DUMMY_10525 AND2_X1 
XU40 CARRYB_15__0_ SUMB_15__1_ n39 NETTRAN_DUMMY_10526 NETTRAN_DUMMY_10527 AND2_X1 
XU39 CARRYB_15__0_ SUMB_15__1_ n38 NETTRAN_DUMMY_10528 NETTRAN_DUMMY_10529 XOR2_X1 
XU38 CARRYB_15__4_ SUMB_15__5_ n37 NETTRAN_DUMMY_10530 NETTRAN_DUMMY_10531 XOR2_X1 
XU37 CARRYB_15__2_ SUMB_15__3_ n36 NETTRAN_DUMMY_10532 NETTRAN_DUMMY_10533 XOR2_X1 
XU36 ab_1__0_ ab_0__1_ PRODUCT[1] NETTRAN_DUMMY_10534 NETTRAN_DUMMY_10535 XOR2_X1 
XU35 CARRYB_15__17_ n70 NETTRAN_DUMMY_10536 NETTRAN_DUMMY_10537 INV_X1 
XU34 ab_1__1_ ab_0__2_ n34 NETTRAN_DUMMY_10538 NETTRAN_DUMMY_10539 XOR2_X1 
XU33 ab_1__2_ ab_0__3_ n33 NETTRAN_DUMMY_10540 NETTRAN_DUMMY_10541 XOR2_X1 
XU32 ab_1__16_ ab_0__17_ n32 NETTRAN_DUMMY_10542 NETTRAN_DUMMY_10543 XOR2_X1 
XU31 ab_1__3_ ab_0__4_ n31 NETTRAN_DUMMY_10544 NETTRAN_DUMMY_10545 XOR2_X1 
XU30 ab_1__4_ ab_0__5_ n30 NETTRAN_DUMMY_10546 NETTRAN_DUMMY_10547 XOR2_X1 
XU29 ab_1__5_ ab_0__6_ n29 NETTRAN_DUMMY_10548 NETTRAN_DUMMY_10549 XOR2_X1 
XU28 ab_1__6_ ab_0__7_ n28 NETTRAN_DUMMY_10550 NETTRAN_DUMMY_10551 XOR2_X1 
XU27 ab_1__7_ ab_0__8_ n27 NETTRAN_DUMMY_10552 NETTRAN_DUMMY_10553 XOR2_X1 
XU26 ab_1__8_ ab_0__9_ n26 NETTRAN_DUMMY_10554 NETTRAN_DUMMY_10555 XOR2_X1 
XU25 ab_1__9_ ab_0__10_ n25 NETTRAN_DUMMY_10556 NETTRAN_DUMMY_10557 XOR2_X1 
XU24 ab_1__10_ ab_0__11_ n24 NETTRAN_DUMMY_10558 NETTRAN_DUMMY_10559 XOR2_X1 
XU23 ab_1__11_ ab_0__12_ n23 NETTRAN_DUMMY_10560 NETTRAN_DUMMY_10561 XOR2_X1 
XU22 ab_1__12_ ab_0__13_ n22 NETTRAN_DUMMY_10562 NETTRAN_DUMMY_10563 XOR2_X1 
XU21 ab_1__13_ ab_0__14_ n21 NETTRAN_DUMMY_10564 NETTRAN_DUMMY_10565 XOR2_X1 
XU20 ab_1__14_ ab_0__15_ n20 NETTRAN_DUMMY_10566 NETTRAN_DUMMY_10567 XOR2_X1 
XU19 ab_1__15_ ab_0__16_ n19 NETTRAN_DUMMY_10568 NETTRAN_DUMMY_10569 XOR2_X1 
XU18 ab_0__17_ ab_1__16_ n18 NETTRAN_DUMMY_10570 NETTRAN_DUMMY_10571 AND2_X1 
XU17 ab_0__1_ ab_1__0_ n17 NETTRAN_DUMMY_10572 NETTRAN_DUMMY_10573 AND2_X1 
XU16 ab_0__2_ ab_1__1_ n16 NETTRAN_DUMMY_10574 NETTRAN_DUMMY_10575 AND2_X1 
XU15 ab_0__3_ ab_1__2_ n15 NETTRAN_DUMMY_10576 NETTRAN_DUMMY_10577 AND2_X1 
XU14 ab_0__4_ ab_1__3_ n14 NETTRAN_DUMMY_10578 NETTRAN_DUMMY_10579 AND2_X1 
XU13 ab_0__5_ ab_1__4_ n13 NETTRAN_DUMMY_10580 NETTRAN_DUMMY_10581 AND2_X1 
XU12 ab_0__6_ ab_1__5_ n12 NETTRAN_DUMMY_10582 NETTRAN_DUMMY_10583 AND2_X1 
XU11 ab_0__7_ ab_1__6_ n11 NETTRAN_DUMMY_10584 NETTRAN_DUMMY_10585 AND2_X1 
XU10 ab_0__8_ ab_1__7_ n10 NETTRAN_DUMMY_10586 NETTRAN_DUMMY_10587 AND2_X1 
XU9 ab_0__9_ ab_1__8_ n9 NETTRAN_DUMMY_10588 NETTRAN_DUMMY_10589 AND2_X1 
XU8 ab_0__10_ ab_1__9_ n8 NETTRAN_DUMMY_10590 NETTRAN_DUMMY_10591 AND2_X1 
XU7 ab_0__11_ ab_1__10_ n7 NETTRAN_DUMMY_10592 NETTRAN_DUMMY_10593 AND2_X1 
XU6 ab_0__12_ ab_1__11_ n6 NETTRAN_DUMMY_10594 NETTRAN_DUMMY_10595 AND2_X1 
XU5 ab_0__13_ ab_1__12_ n5 NETTRAN_DUMMY_10596 NETTRAN_DUMMY_10597 AND2_X1 
XU4 ab_0__14_ ab_1__13_ n4 NETTRAN_DUMMY_10598 NETTRAN_DUMMY_10599 AND2_X1 
XU3 ab_0__15_ ab_1__14_ n3 NETTRAN_DUMMY_10600 NETTRAN_DUMMY_10601 AND2_X1 
XU2 ab_0__16_ ab_1__15_ n2 NETTRAN_DUMMY_10602 NETTRAN_DUMMY_10603 AND2_X1 
XS3_2_16 ab_2__16_ n18 ab_1__17_ CARRYB_2__16_ SUMB_2__16_ NETTRAN_DUMMY_10604 NETTRAN_DUMMY_10605 FA_X1 
XS2_2_15 ab_2__15_ n2 n32 CARRYB_2__15_ SUMB_2__15_ NETTRAN_DUMMY_10606 NETTRAN_DUMMY_10607 FA_X1 
XS2_2_14 ab_2__14_ n3 n19 CARRYB_2__14_ SUMB_2__14_ NETTRAN_DUMMY_10608 NETTRAN_DUMMY_10609 FA_X1 
XS2_2_13 ab_2__13_ n4 n20 CARRYB_2__13_ SUMB_2__13_ NETTRAN_DUMMY_10610 NETTRAN_DUMMY_10611 FA_X1 
XS2_2_12 ab_2__12_ n5 n21 CARRYB_2__12_ SUMB_2__12_ NETTRAN_DUMMY_10612 NETTRAN_DUMMY_10613 FA_X1 
XS2_2_11 ab_2__11_ n6 n22 CARRYB_2__11_ SUMB_2__11_ NETTRAN_DUMMY_10614 NETTRAN_DUMMY_10615 FA_X1 
XS2_2_10 ab_2__10_ n7 n23 CARRYB_2__10_ SUMB_2__10_ NETTRAN_DUMMY_10616 NETTRAN_DUMMY_10617 FA_X1 
XS2_2_9 ab_2__9_ n8 n24 CARRYB_2__9_ SUMB_2__9_ NETTRAN_DUMMY_10618 NETTRAN_DUMMY_10619 FA_X1 
XS2_2_8 ab_2__8_ n9 n25 CARRYB_2__8_ SUMB_2__8_ NETTRAN_DUMMY_10620 NETTRAN_DUMMY_10621 FA_X1 
XS2_2_7 ab_2__7_ n10 n26 CARRYB_2__7_ SUMB_2__7_ NETTRAN_DUMMY_10622 NETTRAN_DUMMY_10623 FA_X1 
XS2_2_6 ab_2__6_ n11 n27 CARRYB_2__6_ SUMB_2__6_ NETTRAN_DUMMY_10624 NETTRAN_DUMMY_10625 FA_X1 
XS2_2_5 ab_2__5_ n12 n28 CARRYB_2__5_ SUMB_2__5_ NETTRAN_DUMMY_10626 NETTRAN_DUMMY_10627 FA_X1 
XS2_2_4 ab_2__4_ n13 n29 CARRYB_2__4_ SUMB_2__4_ NETTRAN_DUMMY_10628 NETTRAN_DUMMY_10629 FA_X1 
XS2_2_3 ab_2__3_ n14 n30 CARRYB_2__3_ SUMB_2__3_ NETTRAN_DUMMY_10630 NETTRAN_DUMMY_10631 FA_X1 
XS2_2_2 ab_2__2_ n15 n31 CARRYB_2__2_ SUMB_2__2_ NETTRAN_DUMMY_10632 NETTRAN_DUMMY_10633 FA_X1 
XS2_2_1 ab_2__1_ n16 n33 CARRYB_2__1_ SUMB_2__1_ NETTRAN_DUMMY_10634 NETTRAN_DUMMY_10635 FA_X1 
XS1_2_0 ab_2__0_ n17 n34 CARRYB_2__0_ PRODUCT[2] NETTRAN_DUMMY_10636 NETTRAN_DUMMY_10637 FA_X1 
XS3_3_16 ab_3__16_ CARRYB_2__16_ ab_2__17_ CARRYB_3__16_ SUMB_3__16_ NETTRAN_DUMMY_10638 
+ NETTRAN_DUMMY_10639 FA_X1 
XS2_3_15 ab_3__15_ CARRYB_2__15_ SUMB_2__16_ CARRYB_3__15_ SUMB_3__15_ NETTRAN_DUMMY_10640 
+ NETTRAN_DUMMY_10641 FA_X1 
XS2_3_14 ab_3__14_ CARRYB_2__14_ SUMB_2__15_ CARRYB_3__14_ SUMB_3__14_ NETTRAN_DUMMY_10642 
+ NETTRAN_DUMMY_10643 FA_X1 
XS2_3_13 ab_3__13_ CARRYB_2__13_ SUMB_2__14_ CARRYB_3__13_ SUMB_3__13_ NETTRAN_DUMMY_10644 
+ NETTRAN_DUMMY_10645 FA_X1 
XS2_3_12 ab_3__12_ CARRYB_2__12_ SUMB_2__13_ CARRYB_3__12_ SUMB_3__12_ NETTRAN_DUMMY_10646 
+ NETTRAN_DUMMY_10647 FA_X1 
XS2_3_11 ab_3__11_ CARRYB_2__11_ SUMB_2__12_ CARRYB_3__11_ SUMB_3__11_ NETTRAN_DUMMY_10648 
+ NETTRAN_DUMMY_10649 FA_X1 
XS2_3_10 ab_3__10_ CARRYB_2__10_ SUMB_2__11_ CARRYB_3__10_ SUMB_3__10_ NETTRAN_DUMMY_10650 
+ NETTRAN_DUMMY_10651 FA_X1 
XS2_3_9 ab_3__9_ CARRYB_2__9_ SUMB_2__10_ CARRYB_3__9_ SUMB_3__9_ NETTRAN_DUMMY_10652 
+ NETTRAN_DUMMY_10653 FA_X1 
XS2_3_8 ab_3__8_ CARRYB_2__8_ SUMB_2__9_ CARRYB_3__8_ SUMB_3__8_ NETTRAN_DUMMY_10654 
+ NETTRAN_DUMMY_10655 FA_X1 
XS2_3_7 ab_3__7_ CARRYB_2__7_ SUMB_2__8_ CARRYB_3__7_ SUMB_3__7_ NETTRAN_DUMMY_10656 
+ NETTRAN_DUMMY_10657 FA_X1 
XS2_3_6 ab_3__6_ CARRYB_2__6_ SUMB_2__7_ CARRYB_3__6_ SUMB_3__6_ NETTRAN_DUMMY_10658 
+ NETTRAN_DUMMY_10659 FA_X1 
XS2_3_5 ab_3__5_ CARRYB_2__5_ SUMB_2__6_ CARRYB_3__5_ SUMB_3__5_ NETTRAN_DUMMY_10660 
+ NETTRAN_DUMMY_10661 FA_X1 
XS2_3_4 ab_3__4_ CARRYB_2__4_ SUMB_2__5_ CARRYB_3__4_ SUMB_3__4_ NETTRAN_DUMMY_10662 
+ NETTRAN_DUMMY_10663 FA_X1 
XS2_3_3 ab_3__3_ CARRYB_2__3_ SUMB_2__4_ CARRYB_3__3_ SUMB_3__3_ NETTRAN_DUMMY_10664 
+ NETTRAN_DUMMY_10665 FA_X1 
XU156 n91 n77 ab_7__11_ NETTRAN_DUMMY_10666 NETTRAN_DUMMY_10667 NOR2_X1 
XU155 n90 n77 ab_7__12_ NETTRAN_DUMMY_10668 NETTRAN_DUMMY_10669 NOR2_X1 
XU154 n89 n77 ab_7__13_ NETTRAN_DUMMY_10670 NETTRAN_DUMMY_10671 NOR2_X1 
XU153 n88 n77 ab_7__14_ NETTRAN_DUMMY_10672 NETTRAN_DUMMY_10673 NOR2_X1 
XU152 n87 n77 ab_7__15_ NETTRAN_DUMMY_10674 NETTRAN_DUMMY_10675 NOR2_X1 
XU151 n86 n77 ab_7__16_ NETTRAN_DUMMY_10676 NETTRAN_DUMMY_10677 NOR2_X1 
XU150 A[7] n85 ab_7__17_ NETTRAN_DUMMY_10678 NETTRAN_DUMMY_10679 NOR2_X1 
XU149 n101 n77 ab_7__1_ NETTRAN_DUMMY_10680 NETTRAN_DUMMY_10681 NOR2_X1 
XU148 n100 n77 ab_7__2_ NETTRAN_DUMMY_10682 NETTRAN_DUMMY_10683 NOR2_X1 
XU147 n99 n77 ab_7__3_ NETTRAN_DUMMY_10684 NETTRAN_DUMMY_10685 NOR2_X1 
XU146 n98 n77 ab_7__4_ NETTRAN_DUMMY_10686 NETTRAN_DUMMY_10687 NOR2_X1 
XU145 n97 n77 ab_7__5_ NETTRAN_DUMMY_10688 NETTRAN_DUMMY_10689 NOR2_X1 
XU144 n96 n77 ab_7__6_ NETTRAN_DUMMY_10690 NETTRAN_DUMMY_10691 NOR2_X1 
XU143 n95 n77 ab_7__7_ NETTRAN_DUMMY_10692 NETTRAN_DUMMY_10693 NOR2_X1 
XU142 n94 n77 ab_7__8_ NETTRAN_DUMMY_10694 NETTRAN_DUMMY_10695 NOR2_X1 
XU141 n93 n77 ab_7__9_ NETTRAN_DUMMY_10696 NETTRAN_DUMMY_10697 NOR2_X1 
XU140 n102 n76 ab_8__0_ NETTRAN_DUMMY_10698 NETTRAN_DUMMY_10699 NOR2_X1 
XU139 n92 n76 ab_8__10_ NETTRAN_DUMMY_10700 NETTRAN_DUMMY_10701 NOR2_X1 
XU138 n91 n76 ab_8__11_ NETTRAN_DUMMY_10702 NETTRAN_DUMMY_10703 NOR2_X1 
XU137 n90 n76 ab_8__12_ NETTRAN_DUMMY_10704 NETTRAN_DUMMY_10705 NOR2_X1 
XU136 n89 n76 ab_8__13_ NETTRAN_DUMMY_10706 NETTRAN_DUMMY_10707 NOR2_X1 
XU135 n88 n76 ab_8__14_ NETTRAN_DUMMY_10708 NETTRAN_DUMMY_10709 NOR2_X1 
XU134 n87 n76 ab_8__15_ NETTRAN_DUMMY_10710 NETTRAN_DUMMY_10711 NOR2_X1 
XU133 n86 n76 ab_8__16_ NETTRAN_DUMMY_10712 NETTRAN_DUMMY_10713 NOR2_X1 
XU132 A[8] n85 ab_8__17_ NETTRAN_DUMMY_10714 NETTRAN_DUMMY_10715 NOR2_X1 
XU131 n101 n76 ab_8__1_ NETTRAN_DUMMY_10716 NETTRAN_DUMMY_10717 NOR2_X1 
XU130 n100 n76 ab_8__2_ NETTRAN_DUMMY_10718 NETTRAN_DUMMY_10719 NOR2_X1 
XU129 n99 n76 ab_8__3_ NETTRAN_DUMMY_10720 NETTRAN_DUMMY_10721 NOR2_X1 
XU128 n98 n76 ab_8__4_ NETTRAN_DUMMY_10722 NETTRAN_DUMMY_10723 NOR2_X1 
XU127 n97 n76 ab_8__5_ NETTRAN_DUMMY_10724 NETTRAN_DUMMY_10725 NOR2_X1 
XU126 n96 n76 ab_8__6_ NETTRAN_DUMMY_10726 NETTRAN_DUMMY_10727 NOR2_X1 
XU125 n95 n76 ab_8__7_ NETTRAN_DUMMY_10728 NETTRAN_DUMMY_10729 NOR2_X1 
XU124 n94 n76 ab_8__8_ NETTRAN_DUMMY_10730 NETTRAN_DUMMY_10731 NOR2_X1 
XU123 n93 n76 ab_8__9_ NETTRAN_DUMMY_10732 NETTRAN_DUMMY_10733 NOR2_X1 
XU122 n75 n102 ab_9__0_ NETTRAN_DUMMY_10734 NETTRAN_DUMMY_10735 NOR2_X1 
XU121 n75 n92 ab_9__10_ NETTRAN_DUMMY_10736 NETTRAN_DUMMY_10737 NOR2_X1 
XU120 n75 n91 ab_9__11_ NETTRAN_DUMMY_10738 NETTRAN_DUMMY_10739 NOR2_X1 
XU119 n75 n90 ab_9__12_ NETTRAN_DUMMY_10740 NETTRAN_DUMMY_10741 NOR2_X1 
XU118 n75 n89 ab_9__13_ NETTRAN_DUMMY_10742 NETTRAN_DUMMY_10743 NOR2_X1 
XU117 n75 n88 ab_9__14_ NETTRAN_DUMMY_10744 NETTRAN_DUMMY_10745 NOR2_X1 
XU116 n75 n87 ab_9__15_ NETTRAN_DUMMY_10746 NETTRAN_DUMMY_10747 NOR2_X1 
XU115 n75 n86 ab_9__16_ NETTRAN_DUMMY_10748 NETTRAN_DUMMY_10749 NOR2_X1 
XU114 A[9] n85 ab_9__17_ NETTRAN_DUMMY_10750 NETTRAN_DUMMY_10751 NOR2_X1 
XU113 n75 n101 ab_9__1_ NETTRAN_DUMMY_10752 NETTRAN_DUMMY_10753 NOR2_X1 
XU112 n75 n100 ab_9__2_ NETTRAN_DUMMY_10754 NETTRAN_DUMMY_10755 NOR2_X1 
XU111 n75 n99 ab_9__3_ NETTRAN_DUMMY_10756 NETTRAN_DUMMY_10757 NOR2_X1 
XU110 n75 n98 ab_9__4_ NETTRAN_DUMMY_10758 NETTRAN_DUMMY_10759 NOR2_X1 
XU109 n75 n97 ab_9__5_ NETTRAN_DUMMY_10760 NETTRAN_DUMMY_10761 NOR2_X1 
XU108 n75 n96 ab_9__6_ NETTRAN_DUMMY_10762 NETTRAN_DUMMY_10763 NOR2_X1 
XU107 n75 n95 ab_9__7_ NETTRAN_DUMMY_10764 NETTRAN_DUMMY_10765 NOR2_X1 
XU106 n75 n94 ab_9__8_ NETTRAN_DUMMY_10766 NETTRAN_DUMMY_10767 NOR2_X1 
XU105 n75 n93 ab_9__9_ NETTRAN_DUMMY_10768 NETTRAN_DUMMY_10769 NOR2_X1 
XU101 A[15] SUMB_15__0_ PRODUCT[15] NETTRAN_DUMMY_10770 NETTRAN_DUMMY_10771 XOR2_X1 
XU89 A[15] SUMB_15__0_ n68 NETTRAN_DUMMY_10772 NETTRAN_DUMMY_10773 AND2_X1 
XU68 CARRYB_15__15_ SUMB_15__16_ n67 NETTRAN_DUMMY_10774 NETTRAN_DUMMY_10775 XOR2_X1 
XU67 CARRYB_15__13_ SUMB_15__14_ n66 NETTRAN_DUMMY_10776 NETTRAN_DUMMY_10777 XOR2_X1 
XU66 CARRYB_15__11_ SUMB_15__12_ n65 NETTRAN_DUMMY_10778 NETTRAN_DUMMY_10779 XOR2_X1 
XU65 CARRYB_15__9_ SUMB_15__10_ n64 NETTRAN_DUMMY_10780 NETTRAN_DUMMY_10781 XOR2_X1 
XU64 CARRYB_15__7_ SUMB_15__8_ n63 NETTRAN_DUMMY_10782 NETTRAN_DUMMY_10783 XOR2_X1 
XU249 n93 n83 ab_1__9_ NETTRAN_DUMMY_10784 NETTRAN_DUMMY_10785 NOR2_X1 
XU248 n102 n82 ab_2__0_ NETTRAN_DUMMY_10786 NETTRAN_DUMMY_10787 NOR2_X1 
XU247 n92 n82 ab_2__10_ NETTRAN_DUMMY_10788 NETTRAN_DUMMY_10789 NOR2_X1 
XU246 n91 n82 ab_2__11_ NETTRAN_DUMMY_10790 NETTRAN_DUMMY_10791 NOR2_X1 
XU245 n90 n82 ab_2__12_ NETTRAN_DUMMY_10792 NETTRAN_DUMMY_10793 NOR2_X1 
XU244 n89 n82 ab_2__13_ NETTRAN_DUMMY_10794 NETTRAN_DUMMY_10795 NOR2_X1 
XU243 n88 n82 ab_2__14_ NETTRAN_DUMMY_10796 NETTRAN_DUMMY_10797 NOR2_X1 
XU242 n87 n82 ab_2__15_ NETTRAN_DUMMY_10798 NETTRAN_DUMMY_10799 NOR2_X1 
XU241 n86 n82 ab_2__16_ NETTRAN_DUMMY_10800 NETTRAN_DUMMY_10801 NOR2_X1 
XU240 A[2] n85 ab_2__17_ NETTRAN_DUMMY_10802 NETTRAN_DUMMY_10803 NOR2_X1 
XU239 n101 n82 ab_2__1_ NETTRAN_DUMMY_10804 NETTRAN_DUMMY_10805 NOR2_X1 
XU238 n100 n82 ab_2__2_ NETTRAN_DUMMY_10806 NETTRAN_DUMMY_10807 NOR2_X1 
XU237 n99 n82 ab_2__3_ NETTRAN_DUMMY_10808 NETTRAN_DUMMY_10809 NOR2_X1 
XU236 n98 n82 ab_2__4_ NETTRAN_DUMMY_10810 NETTRAN_DUMMY_10811 NOR2_X1 
XU235 n97 n82 ab_2__5_ NETTRAN_DUMMY_10812 NETTRAN_DUMMY_10813 NOR2_X1 
XU234 n96 n82 ab_2__6_ NETTRAN_DUMMY_10814 NETTRAN_DUMMY_10815 NOR2_X1 
XU233 n95 n82 ab_2__7_ NETTRAN_DUMMY_10816 NETTRAN_DUMMY_10817 NOR2_X1 
XU232 n94 n82 ab_2__8_ NETTRAN_DUMMY_10818 NETTRAN_DUMMY_10819 NOR2_X1 
XU231 n93 n82 ab_2__9_ NETTRAN_DUMMY_10820 NETTRAN_DUMMY_10821 NOR2_X1 
XU230 n102 n81 ab_3__0_ NETTRAN_DUMMY_10822 NETTRAN_DUMMY_10823 NOR2_X1 
XU229 n92 n81 ab_3__10_ NETTRAN_DUMMY_10824 NETTRAN_DUMMY_10825 NOR2_X1 
XU228 n91 n81 ab_3__11_ NETTRAN_DUMMY_10826 NETTRAN_DUMMY_10827 NOR2_X1 
XU227 n90 n81 ab_3__12_ NETTRAN_DUMMY_10828 NETTRAN_DUMMY_10829 NOR2_X1 
XU226 n89 n81 ab_3__13_ NETTRAN_DUMMY_10830 NETTRAN_DUMMY_10831 NOR2_X1 
XU225 n88 n81 ab_3__14_ NETTRAN_DUMMY_10832 NETTRAN_DUMMY_10833 NOR2_X1 
XU224 n87 n81 ab_3__15_ NETTRAN_DUMMY_10834 NETTRAN_DUMMY_10835 NOR2_X1 
XU223 n86 n81 ab_3__16_ NETTRAN_DUMMY_10836 NETTRAN_DUMMY_10837 NOR2_X1 
XU222 A[3] n85 ab_3__17_ NETTRAN_DUMMY_10838 NETTRAN_DUMMY_10839 NOR2_X1 
XU221 n101 n81 ab_3__1_ NETTRAN_DUMMY_10840 NETTRAN_DUMMY_10841 NOR2_X1 
XU220 n100 n81 ab_3__2_ NETTRAN_DUMMY_10842 NETTRAN_DUMMY_10843 NOR2_X1 
XU219 n99 n81 ab_3__3_ NETTRAN_DUMMY_10844 NETTRAN_DUMMY_10845 NOR2_X1 
XU218 n98 n81 ab_3__4_ NETTRAN_DUMMY_10846 NETTRAN_DUMMY_10847 NOR2_X1 
XU217 n97 n81 ab_3__5_ NETTRAN_DUMMY_10848 NETTRAN_DUMMY_10849 NOR2_X1 
XU216 n96 n81 ab_3__6_ NETTRAN_DUMMY_10850 NETTRAN_DUMMY_10851 NOR2_X1 
XU215 n95 n81 ab_3__7_ NETTRAN_DUMMY_10852 NETTRAN_DUMMY_10853 NOR2_X1 
XU214 n94 n81 ab_3__8_ NETTRAN_DUMMY_10854 NETTRAN_DUMMY_10855 NOR2_X1 
XU213 n93 n81 ab_3__9_ NETTRAN_DUMMY_10856 NETTRAN_DUMMY_10857 NOR2_X1 
XU212 n102 n80 ab_4__0_ NETTRAN_DUMMY_10858 NETTRAN_DUMMY_10859 NOR2_X1 
XU211 n92 n80 ab_4__10_ NETTRAN_DUMMY_10860 NETTRAN_DUMMY_10861 NOR2_X1 
XU210 n91 n80 ab_4__11_ NETTRAN_DUMMY_10862 NETTRAN_DUMMY_10863 NOR2_X1 
XU209 n90 n80 ab_4__12_ NETTRAN_DUMMY_10864 NETTRAN_DUMMY_10865 NOR2_X1 
XU208 n89 n80 ab_4__13_ NETTRAN_DUMMY_10866 NETTRAN_DUMMY_10867 NOR2_X1 
XU207 n88 n80 ab_4__14_ NETTRAN_DUMMY_10868 NETTRAN_DUMMY_10869 NOR2_X1 
XU206 n87 n80 ab_4__15_ NETTRAN_DUMMY_10870 NETTRAN_DUMMY_10871 NOR2_X1 
XU205 n86 n80 ab_4__16_ NETTRAN_DUMMY_10872 NETTRAN_DUMMY_10873 NOR2_X1 
XU204 A[4] n85 ab_4__17_ NETTRAN_DUMMY_10874 NETTRAN_DUMMY_10875 NOR2_X1 
XU203 n101 n80 ab_4__1_ NETTRAN_DUMMY_10876 NETTRAN_DUMMY_10877 NOR2_X1 
XU202 n100 n80 ab_4__2_ NETTRAN_DUMMY_10878 NETTRAN_DUMMY_10879 NOR2_X1 
XU201 n99 n80 ab_4__3_ NETTRAN_DUMMY_10880 NETTRAN_DUMMY_10881 NOR2_X1 
XU200 n98 n80 ab_4__4_ NETTRAN_DUMMY_10882 NETTRAN_DUMMY_10883 NOR2_X1 
XU199 n97 n80 ab_4__5_ NETTRAN_DUMMY_10884 NETTRAN_DUMMY_10885 NOR2_X1 
XU198 n96 n80 ab_4__6_ NETTRAN_DUMMY_10886 NETTRAN_DUMMY_10887 NOR2_X1 
XU197 n95 n80 ab_4__7_ NETTRAN_DUMMY_10888 NETTRAN_DUMMY_10889 NOR2_X1 
XU196 n94 n80 ab_4__8_ NETTRAN_DUMMY_10890 NETTRAN_DUMMY_10891 NOR2_X1 
XU195 n93 n80 ab_4__9_ NETTRAN_DUMMY_10892 NETTRAN_DUMMY_10893 NOR2_X1 
XU194 n102 n79 ab_5__0_ NETTRAN_DUMMY_10894 NETTRAN_DUMMY_10895 NOR2_X1 
XU193 n92 n79 ab_5__10_ NETTRAN_DUMMY_10896 NETTRAN_DUMMY_10897 NOR2_X1 
XU192 n91 n79 ab_5__11_ NETTRAN_DUMMY_10898 NETTRAN_DUMMY_10899 NOR2_X1 
XU191 n90 n79 ab_5__12_ NETTRAN_DUMMY_10900 NETTRAN_DUMMY_10901 NOR2_X1 
XU190 n89 n79 ab_5__13_ NETTRAN_DUMMY_10902 NETTRAN_DUMMY_10903 NOR2_X1 
XU189 n88 n79 ab_5__14_ NETTRAN_DUMMY_10904 NETTRAN_DUMMY_10905 NOR2_X1 
XU188 n87 n79 ab_5__15_ NETTRAN_DUMMY_10906 NETTRAN_DUMMY_10907 NOR2_X1 
XU187 n86 n79 ab_5__16_ NETTRAN_DUMMY_10908 NETTRAN_DUMMY_10909 NOR2_X1 
XU186 A[5] n85 ab_5__17_ NETTRAN_DUMMY_10910 NETTRAN_DUMMY_10911 NOR2_X1 
XU185 n101 n79 ab_5__1_ NETTRAN_DUMMY_10912 NETTRAN_DUMMY_10913 NOR2_X1 
XU184 n100 n79 ab_5__2_ NETTRAN_DUMMY_10914 NETTRAN_DUMMY_10915 NOR2_X1 
XU183 n99 n79 ab_5__3_ NETTRAN_DUMMY_10916 NETTRAN_DUMMY_10917 NOR2_X1 
XU182 n98 n79 ab_5__4_ NETTRAN_DUMMY_10918 NETTRAN_DUMMY_10919 NOR2_X1 
XU181 n97 n79 ab_5__5_ NETTRAN_DUMMY_10920 NETTRAN_DUMMY_10921 NOR2_X1 
XU180 n96 n79 ab_5__6_ NETTRAN_DUMMY_10922 NETTRAN_DUMMY_10923 NOR2_X1 
XU179 n95 n79 ab_5__7_ NETTRAN_DUMMY_10924 NETTRAN_DUMMY_10925 NOR2_X1 
XU178 n94 n79 ab_5__8_ NETTRAN_DUMMY_10926 NETTRAN_DUMMY_10927 NOR2_X1 
XU177 n93 n79 ab_5__9_ NETTRAN_DUMMY_10928 NETTRAN_DUMMY_10929 NOR2_X1 
XU176 n102 n78 ab_6__0_ NETTRAN_DUMMY_10930 NETTRAN_DUMMY_10931 NOR2_X1 
XU175 n92 n78 ab_6__10_ NETTRAN_DUMMY_10932 NETTRAN_DUMMY_10933 NOR2_X1 
XU174 n91 n78 ab_6__11_ NETTRAN_DUMMY_10934 NETTRAN_DUMMY_10935 NOR2_X1 
XU173 n90 n78 ab_6__12_ NETTRAN_DUMMY_10936 NETTRAN_DUMMY_10937 NOR2_X1 
XU172 n89 n78 ab_6__13_ NETTRAN_DUMMY_10938 NETTRAN_DUMMY_10939 NOR2_X1 
XU171 n88 n78 ab_6__14_ NETTRAN_DUMMY_10940 NETTRAN_DUMMY_10941 NOR2_X1 
XU170 n87 n78 ab_6__15_ NETTRAN_DUMMY_10942 NETTRAN_DUMMY_10943 NOR2_X1 
XU169 n86 n78 ab_6__16_ NETTRAN_DUMMY_10944 NETTRAN_DUMMY_10945 NOR2_X1 
XU168 A[6] n85 ab_6__17_ NETTRAN_DUMMY_10946 NETTRAN_DUMMY_10947 NOR2_X1 
XU167 n101 n78 ab_6__1_ NETTRAN_DUMMY_10948 NETTRAN_DUMMY_10949 NOR2_X1 
XU166 n100 n78 ab_6__2_ NETTRAN_DUMMY_10950 NETTRAN_DUMMY_10951 NOR2_X1 
XU165 n99 n78 ab_6__3_ NETTRAN_DUMMY_10952 NETTRAN_DUMMY_10953 NOR2_X1 
XU164 n98 n78 ab_6__4_ NETTRAN_DUMMY_10954 NETTRAN_DUMMY_10955 NOR2_X1 
XU163 n97 n78 ab_6__5_ NETTRAN_DUMMY_10956 NETTRAN_DUMMY_10957 NOR2_X1 
XU162 n96 n78 ab_6__6_ NETTRAN_DUMMY_10958 NETTRAN_DUMMY_10959 NOR2_X1 
XU161 n95 n78 ab_6__7_ NETTRAN_DUMMY_10960 NETTRAN_DUMMY_10961 NOR2_X1 
XU160 n94 n78 ab_6__8_ NETTRAN_DUMMY_10962 NETTRAN_DUMMY_10963 NOR2_X1 
XU159 n93 n78 ab_6__9_ NETTRAN_DUMMY_10964 NETTRAN_DUMMY_10965 NOR2_X1 
XU158 n102 n77 ab_7__0_ NETTRAN_DUMMY_10966 NETTRAN_DUMMY_10967 NOR2_X1 
XU157 n92 n77 ab_7__10_ NETTRAN_DUMMY_10968 NETTRAN_DUMMY_10969 NOR2_X1 
XU342 n96 n73 ab_11__6_ NETTRAN_DUMMY_10970 NETTRAN_DUMMY_10971 NOR2_X1 
XU341 n95 n73 ab_11__7_ NETTRAN_DUMMY_10972 NETTRAN_DUMMY_10973 NOR2_X1 
XU340 n94 n73 ab_11__8_ NETTRAN_DUMMY_10974 NETTRAN_DUMMY_10975 NOR2_X1 
XU339 n93 n73 ab_11__9_ NETTRAN_DUMMY_10976 NETTRAN_DUMMY_10977 NOR2_X1 
XU338 n102 n72 ab_12__0_ NETTRAN_DUMMY_10978 NETTRAN_DUMMY_10979 NOR2_X1 
XU337 n92 n72 ab_12__10_ NETTRAN_DUMMY_10980 NETTRAN_DUMMY_10981 NOR2_X1 
XU336 n91 n72 ab_12__11_ NETTRAN_DUMMY_10982 NETTRAN_DUMMY_10983 NOR2_X1 
XU335 n90 n72 ab_12__12_ NETTRAN_DUMMY_10984 NETTRAN_DUMMY_10985 NOR2_X1 
XU334 n89 n72 ab_12__13_ NETTRAN_DUMMY_10986 NETTRAN_DUMMY_10987 NOR2_X1 
XU333 n88 n72 ab_12__14_ NETTRAN_DUMMY_10988 NETTRAN_DUMMY_10989 NOR2_X1 
XU332 n87 n72 ab_12__15_ NETTRAN_DUMMY_10990 NETTRAN_DUMMY_10991 NOR2_X1 
XU331 n86 n72 ab_12__16_ NETTRAN_DUMMY_10992 NETTRAN_DUMMY_10993 NOR2_X1 
XU330 A[12] n85 ab_12__17_ NETTRAN_DUMMY_10994 NETTRAN_DUMMY_10995 NOR2_X1 
XU329 n101 n72 ab_12__1_ NETTRAN_DUMMY_10996 NETTRAN_DUMMY_10997 NOR2_X1 
XU328 n100 n72 ab_12__2_ NETTRAN_DUMMY_10998 NETTRAN_DUMMY_10999 NOR2_X1 
XU327 n99 n72 ab_12__3_ NETTRAN_DUMMY_11000 NETTRAN_DUMMY_11001 NOR2_X1 
XU326 n98 n72 ab_12__4_ NETTRAN_DUMMY_11002 NETTRAN_DUMMY_11003 NOR2_X1 
XU325 n97 n72 ab_12__5_ NETTRAN_DUMMY_11004 NETTRAN_DUMMY_11005 NOR2_X1 
XU324 n96 n72 ab_12__6_ NETTRAN_DUMMY_11006 NETTRAN_DUMMY_11007 NOR2_X1 
XU323 n95 n72 ab_12__7_ NETTRAN_DUMMY_11008 NETTRAN_DUMMY_11009 NOR2_X1 
XU322 n94 n72 ab_12__8_ NETTRAN_DUMMY_11010 NETTRAN_DUMMY_11011 NOR2_X1 
XU321 n93 n72 ab_12__9_ NETTRAN_DUMMY_11012 NETTRAN_DUMMY_11013 NOR2_X1 
XU320 n102 n71 ab_13__0_ NETTRAN_DUMMY_11014 NETTRAN_DUMMY_11015 NOR2_X1 
XU319 n92 n71 ab_13__10_ NETTRAN_DUMMY_11016 NETTRAN_DUMMY_11017 NOR2_X1 
XU318 n91 n71 ab_13__11_ NETTRAN_DUMMY_11018 NETTRAN_DUMMY_11019 NOR2_X1 
XU317 n90 n71 ab_13__12_ NETTRAN_DUMMY_11020 NETTRAN_DUMMY_11021 NOR2_X1 
XU316 n89 n71 ab_13__13_ NETTRAN_DUMMY_11022 NETTRAN_DUMMY_11023 NOR2_X1 
XU315 n88 n71 ab_13__14_ NETTRAN_DUMMY_11024 NETTRAN_DUMMY_11025 NOR2_X1 
XU314 n87 n71 ab_13__15_ NETTRAN_DUMMY_11026 NETTRAN_DUMMY_11027 NOR2_X1 
XU313 n86 n71 ab_13__16_ NETTRAN_DUMMY_11028 NETTRAN_DUMMY_11029 NOR2_X1 
XU312 A[13] n85 ab_13__17_ NETTRAN_DUMMY_11030 NETTRAN_DUMMY_11031 NOR2_X1 
XU311 n101 n71 ab_13__1_ NETTRAN_DUMMY_11032 NETTRAN_DUMMY_11033 NOR2_X1 
XU310 n100 n71 ab_13__2_ NETTRAN_DUMMY_11034 NETTRAN_DUMMY_11035 NOR2_X1 
XU309 n99 n71 ab_13__3_ NETTRAN_DUMMY_11036 NETTRAN_DUMMY_11037 NOR2_X1 
XU308 n98 n71 ab_13__4_ NETTRAN_DUMMY_11038 NETTRAN_DUMMY_11039 NOR2_X1 
XU307 n97 n71 ab_13__5_ NETTRAN_DUMMY_11040 NETTRAN_DUMMY_11041 NOR2_X1 
XU306 n96 n71 ab_13__6_ NETTRAN_DUMMY_11042 NETTRAN_DUMMY_11043 NOR2_X1 
XU305 n95 n71 ab_13__7_ NETTRAN_DUMMY_11044 NETTRAN_DUMMY_11045 NOR2_X1 
XU304 n94 n71 ab_13__8_ NETTRAN_DUMMY_11046 NETTRAN_DUMMY_11047 NOR2_X1 
XU303 n93 n71 ab_13__9_ NETTRAN_DUMMY_11048 NETTRAN_DUMMY_11049 NOR2_X1 
XU302 n102 n35 ab_14__0_ NETTRAN_DUMMY_11050 NETTRAN_DUMMY_11051 NOR2_X1 
XU301 n92 n35 ab_14__10_ NETTRAN_DUMMY_11052 NETTRAN_DUMMY_11053 NOR2_X1 
XU300 n91 n35 ab_14__11_ NETTRAN_DUMMY_11054 NETTRAN_DUMMY_11055 NOR2_X1 
XU299 n90 n35 ab_14__12_ NETTRAN_DUMMY_11056 NETTRAN_DUMMY_11057 NOR2_X1 
XU298 n89 n35 ab_14__13_ NETTRAN_DUMMY_11058 NETTRAN_DUMMY_11059 NOR2_X1 
XU297 n88 n35 ab_14__14_ NETTRAN_DUMMY_11060 NETTRAN_DUMMY_11061 NOR2_X1 
XU296 n87 n35 ab_14__15_ NETTRAN_DUMMY_11062 NETTRAN_DUMMY_11063 NOR2_X1 
XU295 n86 n35 ab_14__16_ NETTRAN_DUMMY_11064 NETTRAN_DUMMY_11065 NOR2_X1 
XU294 A[14] n85 ab_14__17_ NETTRAN_DUMMY_11066 NETTRAN_DUMMY_11067 NOR2_X1 
XU293 n101 n35 ab_14__1_ NETTRAN_DUMMY_11068 NETTRAN_DUMMY_11069 NOR2_X1 
XU292 n100 n35 ab_14__2_ NETTRAN_DUMMY_11070 NETTRAN_DUMMY_11071 NOR2_X1 
XU291 n99 n35 ab_14__3_ NETTRAN_DUMMY_11072 NETTRAN_DUMMY_11073 NOR2_X1 
XU290 n98 n35 ab_14__4_ NETTRAN_DUMMY_11074 NETTRAN_DUMMY_11075 NOR2_X1 
XU289 n97 n35 ab_14__5_ NETTRAN_DUMMY_11076 NETTRAN_DUMMY_11077 NOR2_X1 
XU288 n96 n35 ab_14__6_ NETTRAN_DUMMY_11078 NETTRAN_DUMMY_11079 NOR2_X1 
XU287 n95 n35 ab_14__7_ NETTRAN_DUMMY_11080 NETTRAN_DUMMY_11081 NOR2_X1 
XU286 n94 n35 ab_14__8_ NETTRAN_DUMMY_11082 NETTRAN_DUMMY_11083 NOR2_X1 
XU285 n93 n35 ab_14__9_ NETTRAN_DUMMY_11084 NETTRAN_DUMMY_11085 NOR2_X1 
XU284 B[0] n1 ab_15__0_ NETTRAN_DUMMY_11086 NETTRAN_DUMMY_11087 NOR2_X1 
XU283 B[10] n1 ab_15__10_ NETTRAN_DUMMY_11088 NETTRAN_DUMMY_11089 NOR2_X1 
XU282 B[11] n1 ab_15__11_ NETTRAN_DUMMY_11090 NETTRAN_DUMMY_11091 NOR2_X1 
XU281 B[12] n1 ab_15__12_ NETTRAN_DUMMY_11092 NETTRAN_DUMMY_11093 NOR2_X1 
XU280 B[13] n1 ab_15__13_ NETTRAN_DUMMY_11094 NETTRAN_DUMMY_11095 NOR2_X1 
XU279 B[14] n1 ab_15__14_ NETTRAN_DUMMY_11096 NETTRAN_DUMMY_11097 NOR2_X1 
XU278 B[15] n1 ab_15__15_ NETTRAN_DUMMY_11098 NETTRAN_DUMMY_11099 NOR2_X1 
XU277 B[16] n1 ab_15__16_ NETTRAN_DUMMY_11100 NETTRAN_DUMMY_11101 NOR2_X1 
XU276 n85 n1 ab_15__17_ NETTRAN_DUMMY_11102 NETTRAN_DUMMY_11103 NOR2_X1 
XU275 B[1] n1 ab_15__1_ NETTRAN_DUMMY_11104 NETTRAN_DUMMY_11105 NOR2_X1 
XU274 B[2] n1 ab_15__2_ NETTRAN_DUMMY_11106 NETTRAN_DUMMY_11107 NOR2_X1 
XU273 B[3] n1 ab_15__3_ NETTRAN_DUMMY_11108 NETTRAN_DUMMY_11109 NOR2_X1 
XU272 B[4] n1 ab_15__4_ NETTRAN_DUMMY_11110 NETTRAN_DUMMY_11111 NOR2_X1 
XU271 B[5] n1 ab_15__5_ NETTRAN_DUMMY_11112 NETTRAN_DUMMY_11113 NOR2_X1 
XU270 B[6] n1 ab_15__6_ NETTRAN_DUMMY_11114 NETTRAN_DUMMY_11115 NOR2_X1 
XU269 B[7] n1 ab_15__7_ NETTRAN_DUMMY_11116 NETTRAN_DUMMY_11117 NOR2_X1 
XU268 B[8] n1 ab_15__8_ NETTRAN_DUMMY_11118 NETTRAN_DUMMY_11119 NOR2_X1 
XU267 B[9] n1 ab_15__9_ NETTRAN_DUMMY_11120 NETTRAN_DUMMY_11121 NOR2_X1 
XU266 n102 n83 ab_1__0_ NETTRAN_DUMMY_11122 NETTRAN_DUMMY_11123 NOR2_X1 
XU265 n92 n83 ab_1__10_ NETTRAN_DUMMY_11124 NETTRAN_DUMMY_11125 NOR2_X1 
XU264 n91 n83 ab_1__11_ NETTRAN_DUMMY_11126 NETTRAN_DUMMY_11127 NOR2_X1 
XU263 n90 n83 ab_1__12_ NETTRAN_DUMMY_11128 NETTRAN_DUMMY_11129 NOR2_X1 
XU262 n89 n83 ab_1__13_ NETTRAN_DUMMY_11130 NETTRAN_DUMMY_11131 NOR2_X1 
XU261 n88 n83 ab_1__14_ NETTRAN_DUMMY_11132 NETTRAN_DUMMY_11133 NOR2_X1 
XU260 n87 n83 ab_1__15_ NETTRAN_DUMMY_11134 NETTRAN_DUMMY_11135 NOR2_X1 
XU259 n86 n83 ab_1__16_ NETTRAN_DUMMY_11136 NETTRAN_DUMMY_11137 NOR2_X1 
XU258 A[1] n85 ab_1__17_ NETTRAN_DUMMY_11138 NETTRAN_DUMMY_11139 NOR2_X1 
XU257 n101 n83 ab_1__1_ NETTRAN_DUMMY_11140 NETTRAN_DUMMY_11141 NOR2_X1 
XU256 n100 n83 ab_1__2_ NETTRAN_DUMMY_11142 NETTRAN_DUMMY_11143 NOR2_X1 
XU255 n99 n83 ab_1__3_ NETTRAN_DUMMY_11144 NETTRAN_DUMMY_11145 NOR2_X1 
XU254 n98 n83 ab_1__4_ NETTRAN_DUMMY_11146 NETTRAN_DUMMY_11147 NOR2_X1 
XU253 n97 n83 ab_1__5_ NETTRAN_DUMMY_11148 NETTRAN_DUMMY_11149 NOR2_X1 
XU252 n96 n83 ab_1__6_ NETTRAN_DUMMY_11150 NETTRAN_DUMMY_11151 NOR2_X1 
XU251 n95 n83 ab_1__7_ NETTRAN_DUMMY_11152 NETTRAN_DUMMY_11153 NOR2_X1 
XU250 n94 n83 ab_1__8_ NETTRAN_DUMMY_11154 NETTRAN_DUMMY_11155 NOR2_X1 
XU392 n102 n84 PRODUCT[0] NETTRAN_DUMMY_11156 NETTRAN_DUMMY_11157 NOR2_X1 
XU391 n92 n84 ab_0__10_ NETTRAN_DUMMY_11158 NETTRAN_DUMMY_11159 NOR2_X1 
XU390 n91 n84 ab_0__11_ NETTRAN_DUMMY_11160 NETTRAN_DUMMY_11161 NOR2_X1 
XU389 n90 n84 ab_0__12_ NETTRAN_DUMMY_11162 NETTRAN_DUMMY_11163 NOR2_X1 
XU388 n89 n84 ab_0__13_ NETTRAN_DUMMY_11164 NETTRAN_DUMMY_11165 NOR2_X1 
XU387 n88 n84 ab_0__14_ NETTRAN_DUMMY_11166 NETTRAN_DUMMY_11167 NOR2_X1 
XU386 n87 n84 ab_0__15_ NETTRAN_DUMMY_11168 NETTRAN_DUMMY_11169 NOR2_X1 
XU385 n86 n84 ab_0__16_ NETTRAN_DUMMY_11170 NETTRAN_DUMMY_11171 NOR2_X1 
XU384 A[0] n85 ab_0__17_ NETTRAN_DUMMY_11172 NETTRAN_DUMMY_11173 NOR2_X1 
XU383 n101 n84 ab_0__1_ NETTRAN_DUMMY_11174 NETTRAN_DUMMY_11175 NOR2_X1 
XU382 n100 n84 ab_0__2_ NETTRAN_DUMMY_11176 NETTRAN_DUMMY_11177 NOR2_X1 
XU381 n99 n84 ab_0__3_ NETTRAN_DUMMY_11178 NETTRAN_DUMMY_11179 NOR2_X1 
XU380 n98 n84 ab_0__4_ NETTRAN_DUMMY_11180 NETTRAN_DUMMY_11181 NOR2_X1 
XU379 n97 n84 ab_0__5_ NETTRAN_DUMMY_11182 NETTRAN_DUMMY_11183 NOR2_X1 
XU378 n96 n84 ab_0__6_ NETTRAN_DUMMY_11184 NETTRAN_DUMMY_11185 NOR2_X1 
XU377 n95 n84 ab_0__7_ NETTRAN_DUMMY_11186 NETTRAN_DUMMY_11187 NOR2_X1 
XU376 n94 n84 ab_0__8_ NETTRAN_DUMMY_11188 NETTRAN_DUMMY_11189 NOR2_X1 
XU375 n93 n84 ab_0__9_ NETTRAN_DUMMY_11190 NETTRAN_DUMMY_11191 NOR2_X1 
XU374 n102 n74 ab_10__0_ NETTRAN_DUMMY_11192 NETTRAN_DUMMY_11193 NOR2_X1 
XU373 n92 n74 ab_10__10_ NETTRAN_DUMMY_11194 NETTRAN_DUMMY_11195 NOR2_X1 
XU372 n91 n74 ab_10__11_ NETTRAN_DUMMY_11196 NETTRAN_DUMMY_11197 NOR2_X1 
XU371 n90 n74 ab_10__12_ NETTRAN_DUMMY_11198 NETTRAN_DUMMY_11199 NOR2_X1 
XU370 n89 n74 ab_10__13_ NETTRAN_DUMMY_11200 NETTRAN_DUMMY_11201 NOR2_X1 
XU369 n88 n74 ab_10__14_ NETTRAN_DUMMY_11202 NETTRAN_DUMMY_11203 NOR2_X1 
XU368 n87 n74 ab_10__15_ NETTRAN_DUMMY_11204 NETTRAN_DUMMY_11205 NOR2_X1 
XU367 n86 n74 ab_10__16_ NETTRAN_DUMMY_11206 NETTRAN_DUMMY_11207 NOR2_X1 
XU366 A[10] n85 ab_10__17_ NETTRAN_DUMMY_11208 NETTRAN_DUMMY_11209 NOR2_X1 
XU365 n101 n74 ab_10__1_ NETTRAN_DUMMY_11210 NETTRAN_DUMMY_11211 NOR2_X1 
XU364 n100 n74 ab_10__2_ NETTRAN_DUMMY_11212 NETTRAN_DUMMY_11213 NOR2_X1 
XU363 n99 n74 ab_10__3_ NETTRAN_DUMMY_11214 NETTRAN_DUMMY_11215 NOR2_X1 
XU362 n98 n74 ab_10__4_ NETTRAN_DUMMY_11216 NETTRAN_DUMMY_11217 NOR2_X1 
XU361 n97 n74 ab_10__5_ NETTRAN_DUMMY_11218 NETTRAN_DUMMY_11219 NOR2_X1 
XU360 n96 n74 ab_10__6_ NETTRAN_DUMMY_11220 NETTRAN_DUMMY_11221 NOR2_X1 
XU359 n95 n74 ab_10__7_ NETTRAN_DUMMY_11222 NETTRAN_DUMMY_11223 NOR2_X1 
XU358 n94 n74 ab_10__8_ NETTRAN_DUMMY_11224 NETTRAN_DUMMY_11225 NOR2_X1 
XU357 n93 n74 ab_10__9_ NETTRAN_DUMMY_11226 NETTRAN_DUMMY_11227 NOR2_X1 
XU356 n102 n73 ab_11__0_ NETTRAN_DUMMY_11228 NETTRAN_DUMMY_11229 NOR2_X1 
XU355 n92 n73 ab_11__10_ NETTRAN_DUMMY_11230 NETTRAN_DUMMY_11231 NOR2_X1 
XU354 n91 n73 ab_11__11_ NETTRAN_DUMMY_11232 NETTRAN_DUMMY_11233 NOR2_X1 
XU353 n90 n73 ab_11__12_ NETTRAN_DUMMY_11234 NETTRAN_DUMMY_11235 NOR2_X1 
XU352 n89 n73 ab_11__13_ NETTRAN_DUMMY_11236 NETTRAN_DUMMY_11237 NOR2_X1 
XU351 n88 n73 ab_11__14_ NETTRAN_DUMMY_11238 NETTRAN_DUMMY_11239 NOR2_X1 
XU350 n87 n73 ab_11__15_ NETTRAN_DUMMY_11240 NETTRAN_DUMMY_11241 NOR2_X1 
XU349 n86 n73 ab_11__16_ NETTRAN_DUMMY_11242 NETTRAN_DUMMY_11243 NOR2_X1 
XU348 A[11] n85 ab_11__17_ NETTRAN_DUMMY_11244 NETTRAN_DUMMY_11245 NOR2_X1 
XU347 n101 n73 ab_11__1_ NETTRAN_DUMMY_11246 NETTRAN_DUMMY_11247 NOR2_X1 
XU346 n100 n73 ab_11__2_ NETTRAN_DUMMY_11248 NETTRAN_DUMMY_11249 NOR2_X1 
XU345 n99 n73 ab_11__3_ NETTRAN_DUMMY_11250 NETTRAN_DUMMY_11251 NOR2_X1 
XU344 n98 n73 ab_11__4_ NETTRAN_DUMMY_11252 NETTRAN_DUMMY_11253 NOR2_X1 
XU343 n97 n73 ab_11__5_ NETTRAN_DUMMY_11254 NETTRAN_DUMMY_11255 NOR2_X1 
XU1 A[15] n1 NETTRAN_DUMMY_11256 NETTRAN_DUMMY_11257 INV_X1 
XU69 A[14] n35 NETTRAN_DUMMY_11258 NETTRAN_DUMMY_11259 INV_X1 
XU70 A[13] n71 NETTRAN_DUMMY_11260 NETTRAN_DUMMY_11261 INV_X1 
XU71 A[12] n72 NETTRAN_DUMMY_11262 NETTRAN_DUMMY_11263 INV_X1 
XU72 A[11] n73 NETTRAN_DUMMY_11264 NETTRAN_DUMMY_11265 INV_X1 
XU73 A[10] n74 NETTRAN_DUMMY_11266 NETTRAN_DUMMY_11267 INV_X1 
XU74 A[9] n75 NETTRAN_DUMMY_11268 NETTRAN_DUMMY_11269 INV_X1 
XU75 A[8] n76 NETTRAN_DUMMY_11270 NETTRAN_DUMMY_11271 INV_X1 
XU76 A[7] n77 NETTRAN_DUMMY_11272 NETTRAN_DUMMY_11273 INV_X1 
XU77 A[6] n78 NETTRAN_DUMMY_11274 NETTRAN_DUMMY_11275 INV_X1 
XU78 A[5] n79 NETTRAN_DUMMY_11276 NETTRAN_DUMMY_11277 INV_X1 
XU79 A[4] n80 NETTRAN_DUMMY_11278 NETTRAN_DUMMY_11279 INV_X1 
XU80 A[3] n81 NETTRAN_DUMMY_11280 NETTRAN_DUMMY_11281 INV_X1 
XU81 A[2] n82 NETTRAN_DUMMY_11282 NETTRAN_DUMMY_11283 INV_X1 
XU82 A[1] n83 NETTRAN_DUMMY_11284 NETTRAN_DUMMY_11285 INV_X1 
XU83 A[0] n84 NETTRAN_DUMMY_11286 NETTRAN_DUMMY_11287 INV_X1 
XU84 B[17] n85 NETTRAN_DUMMY_11288 NETTRAN_DUMMY_11289 INV_X1 
XU85 B[16] n86 NETTRAN_DUMMY_11290 NETTRAN_DUMMY_11291 INV_X1 
XU86 B[15] n87 NETTRAN_DUMMY_11292 NETTRAN_DUMMY_11293 INV_X1 
XU87 B[14] n88 NETTRAN_DUMMY_11294 NETTRAN_DUMMY_11295 INV_X1 
XU88 B[13] n89 NETTRAN_DUMMY_11296 NETTRAN_DUMMY_11297 INV_X1 
XU90 B[12] n90 NETTRAN_DUMMY_11298 NETTRAN_DUMMY_11299 INV_X1 
XU91 B[11] n91 NETTRAN_DUMMY_11300 NETTRAN_DUMMY_11301 INV_X1 
XU92 B[10] n92 NETTRAN_DUMMY_11302 NETTRAN_DUMMY_11303 INV_X1 
XU93 B[9] n93 NETTRAN_DUMMY_11304 NETTRAN_DUMMY_11305 INV_X1 
XU94 B[8] n94 NETTRAN_DUMMY_11306 NETTRAN_DUMMY_11307 INV_X1 
XU95 B[7] n95 NETTRAN_DUMMY_11308 NETTRAN_DUMMY_11309 INV_X1 
XU96 B[6] n96 NETTRAN_DUMMY_11310 NETTRAN_DUMMY_11311 INV_X1 
XU97 B[5] n97 NETTRAN_DUMMY_11312 NETTRAN_DUMMY_11313 INV_X1 
XU98 B[4] n98 NETTRAN_DUMMY_11314 NETTRAN_DUMMY_11315 INV_X1 
XU99 B[3] n99 NETTRAN_DUMMY_11316 NETTRAN_DUMMY_11317 INV_X1 
XU100 B[2] n100 NETTRAN_DUMMY_11318 NETTRAN_DUMMY_11319 INV_X1 
XU102 B[1] n101 NETTRAN_DUMMY_11320 NETTRAN_DUMMY_11321 INV_X1 
XU103 B[0] n102 NETTRAN_DUMMY_11322 NETTRAN_DUMMY_11323 INV_X1 
XFS_1 VSS NETTRAN_DUMMY_11324 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] PRODUCT[29] 
+ PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] PRODUCT[22] 
+ PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] n49 n61 
+ n60 n59 n58 n57 n56 n55 n54 n53 n52 n51 n50 n41 n40 A2_16_ n39 n68 VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS n70 n48 n67 n47 n66 n46 n65 n45 n64 
+ n44 n63 n43 n62 n37 n42 n36 A1_15_ n38 PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] 
+ PRODUCT[11] PRODUCT[10] PRODUCT[9] PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] 
+ PRODUCT[4] PRODUCT[3] PRODUCT[2] gng_smul_16_18_DW01_add_0 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW02_mult_0 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] 
+ PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] PRODUCT[1] 
+ PRODUCT[0] TC B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] 
+ B[5] B[4] B[3] B[2] B[1] B[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] 
+ A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU1 A[15] n1 NETTRAN_DUMMY_11325 NETTRAN_DUMMY_11326 INV_X1 
XS2_11_8 ab_11__8_ CARRYB_10__8_ SUMB_10__9_ CARRYB_11__8_ SUMB_11__8_ NETTRAN_DUMMY_11327 
+ NETTRAN_DUMMY_11328 FA_X1 
XS2_11_7 ab_11__7_ CARRYB_10__7_ SUMB_10__8_ CARRYB_11__7_ SUMB_11__7_ NETTRAN_DUMMY_11329 
+ NETTRAN_DUMMY_11330 FA_X1 
XS2_11_6 ab_11__6_ CARRYB_10__6_ SUMB_10__7_ CARRYB_11__6_ SUMB_11__6_ NETTRAN_DUMMY_11331 
+ NETTRAN_DUMMY_11332 FA_X1 
XS2_11_5 ab_11__5_ CARRYB_10__5_ SUMB_10__6_ CARRYB_11__5_ SUMB_11__5_ NETTRAN_DUMMY_11333 
+ NETTRAN_DUMMY_11334 FA_X1 
XS2_11_4 ab_11__4_ CARRYB_10__4_ SUMB_10__5_ CARRYB_11__4_ SUMB_11__4_ NETTRAN_DUMMY_11335 
+ NETTRAN_DUMMY_11336 FA_X1 
XS2_11_3 ab_11__3_ CARRYB_10__3_ SUMB_10__4_ CARRYB_11__3_ SUMB_11__3_ NETTRAN_DUMMY_11337 
+ NETTRAN_DUMMY_11338 FA_X1 
XS2_11_2 ab_11__2_ CARRYB_10__2_ SUMB_10__3_ CARRYB_11__2_ SUMB_11__2_ NETTRAN_DUMMY_11339 
+ NETTRAN_DUMMY_11340 FA_X1 
XS2_11_1 ab_11__1_ CARRYB_10__1_ SUMB_10__2_ CARRYB_11__1_ SUMB_11__1_ NETTRAN_DUMMY_11341 
+ NETTRAN_DUMMY_11342 FA_X1 
XS1_11_0 ab_11__0_ CARRYB_10__0_ SUMB_10__1_ CARRYB_11__0_ A1_9_ NETTRAN_DUMMY_11343 
+ NETTRAN_DUMMY_11344 FA_X1 
XS3_12_16 ab_12__16_ CARRYB_11__16_ ab_11__17_ CARRYB_12__16_ SUMB_12__16_ NETTRAN_DUMMY_11345 
+ NETTRAN_DUMMY_11346 FA_X1 
XS2_12_15 ab_12__15_ CARRYB_11__15_ SUMB_11__16_ CARRYB_12__15_ SUMB_12__15_ NETTRAN_DUMMY_11347 
+ NETTRAN_DUMMY_11348 FA_X1 
XS2_12_14 ab_12__14_ CARRYB_11__14_ SUMB_11__15_ CARRYB_12__14_ SUMB_12__14_ NETTRAN_DUMMY_11349 
+ NETTRAN_DUMMY_11350 FA_X1 
XS2_12_13 ab_12__13_ CARRYB_11__13_ SUMB_11__14_ CARRYB_12__13_ SUMB_12__13_ NETTRAN_DUMMY_11351 
+ NETTRAN_DUMMY_11352 FA_X1 
XS2_12_12 ab_12__12_ CARRYB_11__12_ SUMB_11__13_ CARRYB_12__12_ SUMB_12__12_ NETTRAN_DUMMY_11353 
+ NETTRAN_DUMMY_11354 FA_X1 
XS2_12_11 ab_12__11_ CARRYB_11__11_ SUMB_11__12_ CARRYB_12__11_ SUMB_12__11_ NETTRAN_DUMMY_11355 
+ NETTRAN_DUMMY_11356 FA_X1 
XS2_12_10 ab_12__10_ CARRYB_11__10_ SUMB_11__11_ CARRYB_12__10_ SUMB_12__10_ NETTRAN_DUMMY_11357 
+ NETTRAN_DUMMY_11358 FA_X1 
XS2_12_9 ab_12__9_ CARRYB_11__9_ SUMB_11__10_ CARRYB_12__9_ SUMB_12__9_ NETTRAN_DUMMY_11359 
+ NETTRAN_DUMMY_11360 FA_X1 
XS2_12_8 ab_12__8_ CARRYB_11__8_ SUMB_11__9_ CARRYB_12__8_ SUMB_12__8_ NETTRAN_DUMMY_11361 
+ NETTRAN_DUMMY_11362 FA_X1 
XS2_12_7 ab_12__7_ CARRYB_11__7_ SUMB_11__8_ CARRYB_12__7_ SUMB_12__7_ NETTRAN_DUMMY_11363 
+ NETTRAN_DUMMY_11364 FA_X1 
XS2_12_6 ab_12__6_ CARRYB_11__6_ SUMB_11__7_ CARRYB_12__6_ SUMB_12__6_ NETTRAN_DUMMY_11365 
+ NETTRAN_DUMMY_11366 FA_X1 
XS2_12_5 ab_12__5_ CARRYB_11__5_ SUMB_11__6_ CARRYB_12__5_ SUMB_12__5_ NETTRAN_DUMMY_11367 
+ NETTRAN_DUMMY_11368 FA_X1 
XS2_12_4 ab_12__4_ CARRYB_11__4_ SUMB_11__5_ CARRYB_12__4_ SUMB_12__4_ NETTRAN_DUMMY_11369 
+ NETTRAN_DUMMY_11370 FA_X1 
XS2_12_3 ab_12__3_ CARRYB_11__3_ SUMB_11__4_ CARRYB_12__3_ SUMB_12__3_ NETTRAN_DUMMY_11371 
+ NETTRAN_DUMMY_11372 FA_X1 
XS2_12_2 ab_12__2_ CARRYB_11__2_ SUMB_11__3_ CARRYB_12__2_ SUMB_12__2_ NETTRAN_DUMMY_11373 
+ NETTRAN_DUMMY_11374 FA_X1 
XS2_12_1 ab_12__1_ CARRYB_11__1_ SUMB_11__2_ CARRYB_12__1_ SUMB_12__1_ NETTRAN_DUMMY_11375 
+ NETTRAN_DUMMY_11376 FA_X1 
XS1_12_0 ab_12__0_ CARRYB_11__0_ SUMB_11__1_ CARRYB_12__0_ A1_10_ NETTRAN_DUMMY_11377 
+ NETTRAN_DUMMY_11378 FA_X1 
XS3_13_16 ab_13__16_ CARRYB_12__16_ ab_12__17_ CARRYB_13__16_ SUMB_13__16_ NETTRAN_DUMMY_11379 
+ NETTRAN_DUMMY_11380 FA_X1 
XS2_13_15 ab_13__15_ CARRYB_12__15_ SUMB_12__16_ CARRYB_13__15_ SUMB_13__15_ NETTRAN_DUMMY_11381 
+ NETTRAN_DUMMY_11382 FA_X1 
XS2_13_14 ab_13__14_ CARRYB_12__14_ SUMB_12__15_ CARRYB_13__14_ SUMB_13__14_ NETTRAN_DUMMY_11383 
+ NETTRAN_DUMMY_11384 FA_X1 
XS2_13_13 ab_13__13_ CARRYB_12__13_ SUMB_12__14_ CARRYB_13__13_ SUMB_13__13_ NETTRAN_DUMMY_11385 
+ NETTRAN_DUMMY_11386 FA_X1 
XS2_13_12 ab_13__12_ CARRYB_12__12_ SUMB_12__13_ CARRYB_13__12_ SUMB_13__12_ NETTRAN_DUMMY_11387 
+ NETTRAN_DUMMY_11388 FA_X1 
XS2_13_11 ab_13__11_ CARRYB_12__11_ SUMB_12__12_ CARRYB_13__11_ SUMB_13__11_ NETTRAN_DUMMY_11389 
+ NETTRAN_DUMMY_11390 FA_X1 
XS2_13_10 ab_13__10_ CARRYB_12__10_ SUMB_12__11_ CARRYB_13__10_ SUMB_13__10_ NETTRAN_DUMMY_11391 
+ NETTRAN_DUMMY_11392 FA_X1 
XS2_13_9 ab_13__9_ CARRYB_12__9_ SUMB_12__10_ CARRYB_13__9_ SUMB_13__9_ NETTRAN_DUMMY_11393 
+ NETTRAN_DUMMY_11394 FA_X1 
XS2_13_8 ab_13__8_ CARRYB_12__8_ SUMB_12__9_ CARRYB_13__8_ SUMB_13__8_ NETTRAN_DUMMY_11395 
+ NETTRAN_DUMMY_11396 FA_X1 
XS2_13_7 ab_13__7_ CARRYB_12__7_ SUMB_12__8_ CARRYB_13__7_ SUMB_13__7_ NETTRAN_DUMMY_11397 
+ NETTRAN_DUMMY_11398 FA_X1 
XS2_13_6 ab_13__6_ CARRYB_12__6_ SUMB_12__7_ CARRYB_13__6_ SUMB_13__6_ NETTRAN_DUMMY_11399 
+ NETTRAN_DUMMY_11400 FA_X1 
XS2_13_5 ab_13__5_ CARRYB_12__5_ SUMB_12__6_ CARRYB_13__5_ SUMB_13__5_ NETTRAN_DUMMY_11401 
+ NETTRAN_DUMMY_11402 FA_X1 
XS2_13_4 ab_13__4_ CARRYB_12__4_ SUMB_12__5_ CARRYB_13__4_ SUMB_13__4_ NETTRAN_DUMMY_11403 
+ NETTRAN_DUMMY_11404 FA_X1 
XS2_13_3 ab_13__3_ CARRYB_12__3_ SUMB_12__4_ CARRYB_13__3_ SUMB_13__3_ NETTRAN_DUMMY_11405 
+ NETTRAN_DUMMY_11406 FA_X1 
XS2_13_2 ab_13__2_ CARRYB_12__2_ SUMB_12__3_ CARRYB_13__2_ SUMB_13__2_ NETTRAN_DUMMY_11407 
+ NETTRAN_DUMMY_11408 FA_X1 
XS2_13_1 ab_13__1_ CARRYB_12__1_ SUMB_12__2_ CARRYB_13__1_ SUMB_13__1_ NETTRAN_DUMMY_11409 
+ NETTRAN_DUMMY_11410 FA_X1 
XS1_13_0 ab_13__0_ CARRYB_12__0_ SUMB_12__1_ CARRYB_13__0_ A1_11_ NETTRAN_DUMMY_11411 
+ NETTRAN_DUMMY_11412 FA_X1 
XS3_14_16 ab_14__16_ CARRYB_13__16_ ab_13__17_ CARRYB_14__16_ SUMB_14__16_ NETTRAN_DUMMY_11413 
+ NETTRAN_DUMMY_11414 FA_X1 
XS2_14_15 ab_14__15_ CARRYB_13__15_ SUMB_13__16_ CARRYB_14__15_ SUMB_14__15_ NETTRAN_DUMMY_11415 
+ NETTRAN_DUMMY_11416 FA_X1 
XS2_14_14 ab_14__14_ CARRYB_13__14_ SUMB_13__15_ CARRYB_14__14_ SUMB_14__14_ NETTRAN_DUMMY_11417 
+ NETTRAN_DUMMY_11418 FA_X1 
XS2_14_13 ab_14__13_ CARRYB_13__13_ SUMB_13__14_ CARRYB_14__13_ SUMB_14__13_ NETTRAN_DUMMY_11419 
+ NETTRAN_DUMMY_11420 FA_X1 
XS2_14_12 ab_14__12_ CARRYB_13__12_ SUMB_13__13_ CARRYB_14__12_ SUMB_14__12_ NETTRAN_DUMMY_11421 
+ NETTRAN_DUMMY_11422 FA_X1 
XS2_14_11 ab_14__11_ CARRYB_13__11_ SUMB_13__12_ CARRYB_14__11_ SUMB_14__11_ NETTRAN_DUMMY_11423 
+ NETTRAN_DUMMY_11424 FA_X1 
XS2_14_10 ab_14__10_ CARRYB_13__10_ SUMB_13__11_ CARRYB_14__10_ SUMB_14__10_ NETTRAN_DUMMY_11425 
+ NETTRAN_DUMMY_11426 FA_X1 
XS2_14_9 ab_14__9_ CARRYB_13__9_ SUMB_13__10_ CARRYB_14__9_ SUMB_14__9_ NETTRAN_DUMMY_11427 
+ NETTRAN_DUMMY_11428 FA_X1 
XS2_14_8 ab_14__8_ CARRYB_13__8_ SUMB_13__9_ CARRYB_14__8_ SUMB_14__8_ NETTRAN_DUMMY_11429 
+ NETTRAN_DUMMY_11430 FA_X1 
XS2_14_7 ab_14__7_ CARRYB_13__7_ SUMB_13__8_ CARRYB_14__7_ SUMB_14__7_ NETTRAN_DUMMY_11431 
+ NETTRAN_DUMMY_11432 FA_X1 
XS2_14_6 ab_14__6_ CARRYB_13__6_ SUMB_13__7_ CARRYB_14__6_ SUMB_14__6_ NETTRAN_DUMMY_11433 
+ NETTRAN_DUMMY_11434 FA_X1 
XS2_14_5 ab_14__5_ CARRYB_13__5_ SUMB_13__6_ CARRYB_14__5_ SUMB_14__5_ NETTRAN_DUMMY_11435 
+ NETTRAN_DUMMY_11436 FA_X1 
XS2_14_4 ab_14__4_ CARRYB_13__4_ SUMB_13__5_ CARRYB_14__4_ SUMB_14__4_ NETTRAN_DUMMY_11437 
+ NETTRAN_DUMMY_11438 FA_X1 
XS2_14_3 ab_14__3_ CARRYB_13__3_ SUMB_13__4_ CARRYB_14__3_ SUMB_14__3_ NETTRAN_DUMMY_11439 
+ NETTRAN_DUMMY_11440 FA_X1 
XS2_14_2 ab_14__2_ CARRYB_13__2_ SUMB_13__3_ CARRYB_14__2_ SUMB_14__2_ NETTRAN_DUMMY_11441 
+ NETTRAN_DUMMY_11442 FA_X1 
XS2_14_1 ab_14__1_ CARRYB_13__1_ SUMB_13__2_ CARRYB_14__1_ SUMB_14__1_ NETTRAN_DUMMY_11443 
+ NETTRAN_DUMMY_11444 FA_X1 
XS1_14_0 ab_14__0_ CARRYB_13__0_ SUMB_13__1_ CARRYB_14__0_ A1_12_ NETTRAN_DUMMY_11445 
+ NETTRAN_DUMMY_11446 FA_X1 
XS14_17 n1 n85 ab_15__17_ CARRYB_15__17_ SUMB_15__17_ NETTRAN_DUMMY_11447 NETTRAN_DUMMY_11448 FA_X1 
XS5_16 ab_15__16_ CARRYB_14__16_ ab_14__17_ CARRYB_15__16_ SUMB_15__16_ NETTRAN_DUMMY_11449 
+ NETTRAN_DUMMY_11450 FA_X1 
XS4_15 ab_15__15_ CARRYB_14__15_ SUMB_14__16_ CARRYB_15__15_ SUMB_15__15_ NETTRAN_DUMMY_11451 
+ NETTRAN_DUMMY_11452 FA_X1 
XS4_14 ab_15__14_ CARRYB_14__14_ SUMB_14__15_ CARRYB_15__14_ SUMB_15__14_ NETTRAN_DUMMY_11453 
+ NETTRAN_DUMMY_11454 FA_X1 
XS4_13 ab_15__13_ CARRYB_14__13_ SUMB_14__14_ CARRYB_15__13_ SUMB_15__13_ NETTRAN_DUMMY_11455 
+ NETTRAN_DUMMY_11456 FA_X1 
XS4_12 ab_15__12_ CARRYB_14__12_ SUMB_14__13_ CARRYB_15__12_ SUMB_15__12_ NETTRAN_DUMMY_11457 
+ NETTRAN_DUMMY_11458 FA_X1 
XS4_11 ab_15__11_ CARRYB_14__11_ SUMB_14__12_ CARRYB_15__11_ SUMB_15__11_ NETTRAN_DUMMY_11459 
+ NETTRAN_DUMMY_11460 FA_X1 
XS4_10 ab_15__10_ CARRYB_14__10_ SUMB_14__11_ CARRYB_15__10_ SUMB_15__10_ NETTRAN_DUMMY_11461 
+ NETTRAN_DUMMY_11462 FA_X1 
XS4_9 ab_15__9_ CARRYB_14__9_ SUMB_14__10_ CARRYB_15__9_ SUMB_15__9_ NETTRAN_DUMMY_11463 
+ NETTRAN_DUMMY_11464 FA_X1 
XS4_8 ab_15__8_ CARRYB_14__8_ SUMB_14__9_ CARRYB_15__8_ SUMB_15__8_ NETTRAN_DUMMY_11465 
+ NETTRAN_DUMMY_11466 FA_X1 
XS4_7 ab_15__7_ CARRYB_14__7_ SUMB_14__8_ CARRYB_15__7_ SUMB_15__7_ NETTRAN_DUMMY_11467 
+ NETTRAN_DUMMY_11468 FA_X1 
XS4_6 ab_15__6_ CARRYB_14__6_ SUMB_14__7_ CARRYB_15__6_ SUMB_15__6_ NETTRAN_DUMMY_11469 
+ NETTRAN_DUMMY_11470 FA_X1 
XS4_5 ab_15__5_ CARRYB_14__5_ SUMB_14__6_ CARRYB_15__5_ SUMB_15__5_ NETTRAN_DUMMY_11471 
+ NETTRAN_DUMMY_11472 FA_X1 
XS4_4 ab_15__4_ CARRYB_14__4_ SUMB_14__5_ CARRYB_15__4_ SUMB_15__4_ NETTRAN_DUMMY_11473 
+ NETTRAN_DUMMY_11474 FA_X1 
XS4_3 ab_15__3_ CARRYB_14__3_ SUMB_14__4_ CARRYB_15__3_ SUMB_15__3_ NETTRAN_DUMMY_11475 
+ NETTRAN_DUMMY_11476 FA_X1 
XS4_2 ab_15__2_ CARRYB_14__2_ SUMB_14__3_ CARRYB_15__2_ SUMB_15__2_ NETTRAN_DUMMY_11477 
+ NETTRAN_DUMMY_11478 FA_X1 
XS4_1 ab_15__1_ CARRYB_14__1_ SUMB_14__2_ CARRYB_15__1_ SUMB_15__1_ NETTRAN_DUMMY_11479 
+ NETTRAN_DUMMY_11480 FA_X1 
XS4_0 ab_15__0_ CARRYB_14__0_ SUMB_14__1_ CARRYB_15__0_ SUMB_15__0_ NETTRAN_DUMMY_11481 
+ NETTRAN_DUMMY_11482 FA_X1 
XS14_17_0 B[17] CARRYB_15__1_ SUMB_15__2_ A2_16_ A1_15_ NETTRAN_DUMMY_11483 NETTRAN_DUMMY_11484 FA_X1 
XS3_6_16 ab_6__16_ CARRYB_5__16_ ab_5__17_ CARRYB_6__16_ SUMB_6__16_ NETTRAN_DUMMY_11485 
+ NETTRAN_DUMMY_11486 FA_X1 
XS2_6_15 ab_6__15_ CARRYB_5__15_ SUMB_5__16_ CARRYB_6__15_ SUMB_6__15_ NETTRAN_DUMMY_11487 
+ NETTRAN_DUMMY_11488 FA_X1 
XS2_6_14 ab_6__14_ CARRYB_5__14_ SUMB_5__15_ CARRYB_6__14_ SUMB_6__14_ NETTRAN_DUMMY_11489 
+ NETTRAN_DUMMY_11490 FA_X1 
XS2_6_13 ab_6__13_ CARRYB_5__13_ SUMB_5__14_ CARRYB_6__13_ SUMB_6__13_ NETTRAN_DUMMY_11491 
+ NETTRAN_DUMMY_11492 FA_X1 
XS2_6_12 ab_6__12_ CARRYB_5__12_ SUMB_5__13_ CARRYB_6__12_ SUMB_6__12_ NETTRAN_DUMMY_11493 
+ NETTRAN_DUMMY_11494 FA_X1 
XS2_6_11 ab_6__11_ CARRYB_5__11_ SUMB_5__12_ CARRYB_6__11_ SUMB_6__11_ NETTRAN_DUMMY_11495 
+ NETTRAN_DUMMY_11496 FA_X1 
XS2_6_10 ab_6__10_ CARRYB_5__10_ SUMB_5__11_ CARRYB_6__10_ SUMB_6__10_ NETTRAN_DUMMY_11497 
+ NETTRAN_DUMMY_11498 FA_X1 
XS2_6_9 ab_6__9_ CARRYB_5__9_ SUMB_5__10_ CARRYB_6__9_ SUMB_6__9_ NETTRAN_DUMMY_11499 
+ NETTRAN_DUMMY_11500 FA_X1 
XS2_6_8 ab_6__8_ CARRYB_5__8_ SUMB_5__9_ CARRYB_6__8_ SUMB_6__8_ NETTRAN_DUMMY_11501 
+ NETTRAN_DUMMY_11502 FA_X1 
XS2_6_7 ab_6__7_ CARRYB_5__7_ SUMB_5__8_ CARRYB_6__7_ SUMB_6__7_ NETTRAN_DUMMY_11503 
+ NETTRAN_DUMMY_11504 FA_X1 
XS2_6_6 ab_6__6_ CARRYB_5__6_ SUMB_5__7_ CARRYB_6__6_ SUMB_6__6_ NETTRAN_DUMMY_11505 
+ NETTRAN_DUMMY_11506 FA_X1 
XS2_6_5 ab_6__5_ CARRYB_5__5_ SUMB_5__6_ CARRYB_6__5_ SUMB_6__5_ NETTRAN_DUMMY_11507 
+ NETTRAN_DUMMY_11508 FA_X1 
XS2_6_4 ab_6__4_ CARRYB_5__4_ SUMB_5__5_ CARRYB_6__4_ SUMB_6__4_ NETTRAN_DUMMY_11509 
+ NETTRAN_DUMMY_11510 FA_X1 
XS2_6_3 ab_6__3_ CARRYB_5__3_ SUMB_5__4_ CARRYB_6__3_ SUMB_6__3_ NETTRAN_DUMMY_11511 
+ NETTRAN_DUMMY_11512 FA_X1 
XS2_6_2 ab_6__2_ CARRYB_5__2_ SUMB_5__3_ CARRYB_6__2_ SUMB_6__2_ NETTRAN_DUMMY_11513 
+ NETTRAN_DUMMY_11514 FA_X1 
XS2_6_1 ab_6__1_ CARRYB_5__1_ SUMB_5__2_ CARRYB_6__1_ SUMB_6__1_ NETTRAN_DUMMY_11515 
+ NETTRAN_DUMMY_11516 FA_X1 
XS1_6_0 ab_6__0_ CARRYB_5__0_ SUMB_5__1_ CARRYB_6__0_ A1_4_ NETTRAN_DUMMY_11517 
+ NETTRAN_DUMMY_11518 FA_X1 
XS3_7_16 ab_7__16_ CARRYB_6__16_ ab_6__17_ CARRYB_7__16_ SUMB_7__16_ NETTRAN_DUMMY_11519 
+ NETTRAN_DUMMY_11520 FA_X1 
XS2_7_15 ab_7__15_ CARRYB_6__15_ SUMB_6__16_ CARRYB_7__15_ SUMB_7__15_ NETTRAN_DUMMY_11521 
+ NETTRAN_DUMMY_11522 FA_X1 
XS2_7_14 ab_7__14_ CARRYB_6__14_ SUMB_6__15_ CARRYB_7__14_ SUMB_7__14_ NETTRAN_DUMMY_11523 
+ NETTRAN_DUMMY_11524 FA_X1 
XS2_7_13 ab_7__13_ CARRYB_6__13_ SUMB_6__14_ CARRYB_7__13_ SUMB_7__13_ NETTRAN_DUMMY_11525 
+ NETTRAN_DUMMY_11526 FA_X1 
XS2_7_12 ab_7__12_ CARRYB_6__12_ SUMB_6__13_ CARRYB_7__12_ SUMB_7__12_ NETTRAN_DUMMY_11527 
+ NETTRAN_DUMMY_11528 FA_X1 
XS2_7_11 ab_7__11_ CARRYB_6__11_ SUMB_6__12_ CARRYB_7__11_ SUMB_7__11_ NETTRAN_DUMMY_11529 
+ NETTRAN_DUMMY_11530 FA_X1 
XS2_7_10 ab_7__10_ CARRYB_6__10_ SUMB_6__11_ CARRYB_7__10_ SUMB_7__10_ NETTRAN_DUMMY_11531 
+ NETTRAN_DUMMY_11532 FA_X1 
XS2_7_9 ab_7__9_ CARRYB_6__9_ SUMB_6__10_ CARRYB_7__9_ SUMB_7__9_ NETTRAN_DUMMY_11533 
+ NETTRAN_DUMMY_11534 FA_X1 
XS2_7_8 ab_7__8_ CARRYB_6__8_ SUMB_6__9_ CARRYB_7__8_ SUMB_7__8_ NETTRAN_DUMMY_11535 
+ NETTRAN_DUMMY_11536 FA_X1 
XS2_7_7 ab_7__7_ CARRYB_6__7_ SUMB_6__8_ CARRYB_7__7_ SUMB_7__7_ NETTRAN_DUMMY_11537 
+ NETTRAN_DUMMY_11538 FA_X1 
XS2_7_6 ab_7__6_ CARRYB_6__6_ SUMB_6__7_ CARRYB_7__6_ SUMB_7__6_ NETTRAN_DUMMY_11539 
+ NETTRAN_DUMMY_11540 FA_X1 
XS2_7_5 ab_7__5_ CARRYB_6__5_ SUMB_6__6_ CARRYB_7__5_ SUMB_7__5_ NETTRAN_DUMMY_11541 
+ NETTRAN_DUMMY_11542 FA_X1 
XS2_7_4 ab_7__4_ CARRYB_6__4_ SUMB_6__5_ CARRYB_7__4_ SUMB_7__4_ NETTRAN_DUMMY_11543 
+ NETTRAN_DUMMY_11544 FA_X1 
XS2_7_3 ab_7__3_ CARRYB_6__3_ SUMB_6__4_ CARRYB_7__3_ SUMB_7__3_ NETTRAN_DUMMY_11545 
+ NETTRAN_DUMMY_11546 FA_X1 
XS2_7_2 ab_7__2_ CARRYB_6__2_ SUMB_6__3_ CARRYB_7__2_ SUMB_7__2_ NETTRAN_DUMMY_11547 
+ NETTRAN_DUMMY_11548 FA_X1 
XS2_7_1 ab_7__1_ CARRYB_6__1_ SUMB_6__2_ CARRYB_7__1_ SUMB_7__1_ NETTRAN_DUMMY_11549 
+ NETTRAN_DUMMY_11550 FA_X1 
XS1_7_0 ab_7__0_ CARRYB_6__0_ SUMB_6__1_ CARRYB_7__0_ A1_5_ NETTRAN_DUMMY_11551 
+ NETTRAN_DUMMY_11552 FA_X1 
XS3_8_16 ab_8__16_ CARRYB_7__16_ ab_7__17_ CARRYB_8__16_ SUMB_8__16_ NETTRAN_DUMMY_11553 
+ NETTRAN_DUMMY_11554 FA_X1 
XS2_8_15 ab_8__15_ CARRYB_7__15_ SUMB_7__16_ CARRYB_8__15_ SUMB_8__15_ NETTRAN_DUMMY_11555 
+ NETTRAN_DUMMY_11556 FA_X1 
XS2_8_14 ab_8__14_ CARRYB_7__14_ SUMB_7__15_ CARRYB_8__14_ SUMB_8__14_ NETTRAN_DUMMY_11557 
+ NETTRAN_DUMMY_11558 FA_X1 
XS2_8_13 ab_8__13_ CARRYB_7__13_ SUMB_7__14_ CARRYB_8__13_ SUMB_8__13_ NETTRAN_DUMMY_11559 
+ NETTRAN_DUMMY_11560 FA_X1 
XS2_8_12 ab_8__12_ CARRYB_7__12_ SUMB_7__13_ CARRYB_8__12_ SUMB_8__12_ NETTRAN_DUMMY_11561 
+ NETTRAN_DUMMY_11562 FA_X1 
XS2_8_11 ab_8__11_ CARRYB_7__11_ SUMB_7__12_ CARRYB_8__11_ SUMB_8__11_ NETTRAN_DUMMY_11563 
+ NETTRAN_DUMMY_11564 FA_X1 
XS2_8_10 ab_8__10_ CARRYB_7__10_ SUMB_7__11_ CARRYB_8__10_ SUMB_8__10_ NETTRAN_DUMMY_11565 
+ NETTRAN_DUMMY_11566 FA_X1 
XS2_8_9 ab_8__9_ CARRYB_7__9_ SUMB_7__10_ CARRYB_8__9_ SUMB_8__9_ NETTRAN_DUMMY_11567 
+ NETTRAN_DUMMY_11568 FA_X1 
XS2_8_8 ab_8__8_ CARRYB_7__8_ SUMB_7__9_ CARRYB_8__8_ SUMB_8__8_ NETTRAN_DUMMY_11569 
+ NETTRAN_DUMMY_11570 FA_X1 
XS2_8_7 ab_8__7_ CARRYB_7__7_ SUMB_7__8_ CARRYB_8__7_ SUMB_8__7_ NETTRAN_DUMMY_11571 
+ NETTRAN_DUMMY_11572 FA_X1 
XS2_8_6 ab_8__6_ CARRYB_7__6_ SUMB_7__7_ CARRYB_8__6_ SUMB_8__6_ NETTRAN_DUMMY_11573 
+ NETTRAN_DUMMY_11574 FA_X1 
XS2_8_5 ab_8__5_ CARRYB_7__5_ SUMB_7__6_ CARRYB_8__5_ SUMB_8__5_ NETTRAN_DUMMY_11575 
+ NETTRAN_DUMMY_11576 FA_X1 
XS2_8_4 ab_8__4_ CARRYB_7__4_ SUMB_7__5_ CARRYB_8__4_ SUMB_8__4_ NETTRAN_DUMMY_11577 
+ NETTRAN_DUMMY_11578 FA_X1 
XS2_8_3 ab_8__3_ CARRYB_7__3_ SUMB_7__4_ CARRYB_8__3_ SUMB_8__3_ NETTRAN_DUMMY_11579 
+ NETTRAN_DUMMY_11580 FA_X1 
XS2_8_2 ab_8__2_ CARRYB_7__2_ SUMB_7__3_ CARRYB_8__2_ SUMB_8__2_ NETTRAN_DUMMY_11581 
+ NETTRAN_DUMMY_11582 FA_X1 
XS2_8_1 ab_8__1_ CARRYB_7__1_ SUMB_7__2_ CARRYB_8__1_ SUMB_8__1_ NETTRAN_DUMMY_11583 
+ NETTRAN_DUMMY_11584 FA_X1 
XS1_8_0 ab_8__0_ CARRYB_7__0_ SUMB_7__1_ CARRYB_8__0_ A1_6_ NETTRAN_DUMMY_11585 
+ NETTRAN_DUMMY_11586 FA_X1 
XS3_9_16 ab_9__16_ CARRYB_8__16_ ab_8__17_ CARRYB_9__16_ SUMB_9__16_ NETTRAN_DUMMY_11587 
+ NETTRAN_DUMMY_11588 FA_X1 
XS2_9_15 ab_9__15_ CARRYB_8__15_ SUMB_8__16_ CARRYB_9__15_ SUMB_9__15_ NETTRAN_DUMMY_11589 
+ NETTRAN_DUMMY_11590 FA_X1 
XS2_9_14 ab_9__14_ CARRYB_8__14_ SUMB_8__15_ CARRYB_9__14_ SUMB_9__14_ NETTRAN_DUMMY_11591 
+ NETTRAN_DUMMY_11592 FA_X1 
XS2_9_13 ab_9__13_ CARRYB_8__13_ SUMB_8__14_ CARRYB_9__13_ SUMB_9__13_ NETTRAN_DUMMY_11593 
+ NETTRAN_DUMMY_11594 FA_X1 
XS2_9_12 ab_9__12_ CARRYB_8__12_ SUMB_8__13_ CARRYB_9__12_ SUMB_9__12_ NETTRAN_DUMMY_11595 
+ NETTRAN_DUMMY_11596 FA_X1 
XS2_9_11 ab_9__11_ CARRYB_8__11_ SUMB_8__12_ CARRYB_9__11_ SUMB_9__11_ NETTRAN_DUMMY_11597 
+ NETTRAN_DUMMY_11598 FA_X1 
XS2_9_10 ab_9__10_ CARRYB_8__10_ SUMB_8__11_ CARRYB_9__10_ SUMB_9__10_ NETTRAN_DUMMY_11599 
+ NETTRAN_DUMMY_11600 FA_X1 
XS2_9_9 ab_9__9_ CARRYB_8__9_ SUMB_8__10_ CARRYB_9__9_ SUMB_9__9_ NETTRAN_DUMMY_11601 
+ NETTRAN_DUMMY_11602 FA_X1 
XS2_9_8 ab_9__8_ CARRYB_8__8_ SUMB_8__9_ CARRYB_9__8_ SUMB_9__8_ NETTRAN_DUMMY_11603 
+ NETTRAN_DUMMY_11604 FA_X1 
XS2_9_7 ab_9__7_ CARRYB_8__7_ SUMB_8__8_ CARRYB_9__7_ SUMB_9__7_ NETTRAN_DUMMY_11605 
+ NETTRAN_DUMMY_11606 FA_X1 
XS2_9_6 ab_9__6_ CARRYB_8__6_ SUMB_8__7_ CARRYB_9__6_ SUMB_9__6_ NETTRAN_DUMMY_11607 
+ NETTRAN_DUMMY_11608 FA_X1 
XS2_9_5 ab_9__5_ CARRYB_8__5_ SUMB_8__6_ CARRYB_9__5_ SUMB_9__5_ NETTRAN_DUMMY_11609 
+ NETTRAN_DUMMY_11610 FA_X1 
XS2_9_4 ab_9__4_ CARRYB_8__4_ SUMB_8__5_ CARRYB_9__4_ SUMB_9__4_ NETTRAN_DUMMY_11611 
+ NETTRAN_DUMMY_11612 FA_X1 
XS2_9_3 ab_9__3_ CARRYB_8__3_ SUMB_8__4_ CARRYB_9__3_ SUMB_9__3_ NETTRAN_DUMMY_11613 
+ NETTRAN_DUMMY_11614 FA_X1 
XS2_9_2 ab_9__2_ CARRYB_8__2_ SUMB_8__3_ CARRYB_9__2_ SUMB_9__2_ NETTRAN_DUMMY_11615 
+ NETTRAN_DUMMY_11616 FA_X1 
XS2_9_1 ab_9__1_ CARRYB_8__1_ SUMB_8__2_ CARRYB_9__1_ SUMB_9__1_ NETTRAN_DUMMY_11617 
+ NETTRAN_DUMMY_11618 FA_X1 
XS1_9_0 ab_9__0_ CARRYB_8__0_ SUMB_8__1_ CARRYB_9__0_ A1_7_ NETTRAN_DUMMY_11619 
+ NETTRAN_DUMMY_11620 FA_X1 
XS3_10_16 ab_10__16_ CARRYB_9__16_ ab_9__17_ CARRYB_10__16_ SUMB_10__16_ NETTRAN_DUMMY_11621 
+ NETTRAN_DUMMY_11622 FA_X1 
XS2_10_15 ab_10__15_ CARRYB_9__15_ SUMB_9__16_ CARRYB_10__15_ SUMB_10__15_ NETTRAN_DUMMY_11623 
+ NETTRAN_DUMMY_11624 FA_X1 
XS2_10_14 ab_10__14_ CARRYB_9__14_ SUMB_9__15_ CARRYB_10__14_ SUMB_10__14_ NETTRAN_DUMMY_11625 
+ NETTRAN_DUMMY_11626 FA_X1 
XS2_10_13 ab_10__13_ CARRYB_9__13_ SUMB_9__14_ CARRYB_10__13_ SUMB_10__13_ NETTRAN_DUMMY_11627 
+ NETTRAN_DUMMY_11628 FA_X1 
XS2_10_12 ab_10__12_ CARRYB_9__12_ SUMB_9__13_ CARRYB_10__12_ SUMB_10__12_ NETTRAN_DUMMY_11629 
+ NETTRAN_DUMMY_11630 FA_X1 
XS2_10_11 ab_10__11_ CARRYB_9__11_ SUMB_9__12_ CARRYB_10__11_ SUMB_10__11_ NETTRAN_DUMMY_11631 
+ NETTRAN_DUMMY_11632 FA_X1 
XS2_10_10 ab_10__10_ CARRYB_9__10_ SUMB_9__11_ CARRYB_10__10_ SUMB_10__10_ NETTRAN_DUMMY_11633 
+ NETTRAN_DUMMY_11634 FA_X1 
XS2_10_9 ab_10__9_ CARRYB_9__9_ SUMB_9__10_ CARRYB_10__9_ SUMB_10__9_ NETTRAN_DUMMY_11635 
+ NETTRAN_DUMMY_11636 FA_X1 
XS2_10_8 ab_10__8_ CARRYB_9__8_ SUMB_9__9_ CARRYB_10__8_ SUMB_10__8_ NETTRAN_DUMMY_11637 
+ NETTRAN_DUMMY_11638 FA_X1 
XS2_10_7 ab_10__7_ CARRYB_9__7_ SUMB_9__8_ CARRYB_10__7_ SUMB_10__7_ NETTRAN_DUMMY_11639 
+ NETTRAN_DUMMY_11640 FA_X1 
XS2_10_6 ab_10__6_ CARRYB_9__6_ SUMB_9__7_ CARRYB_10__6_ SUMB_10__6_ NETTRAN_DUMMY_11641 
+ NETTRAN_DUMMY_11642 FA_X1 
XS2_10_5 ab_10__5_ CARRYB_9__5_ SUMB_9__6_ CARRYB_10__5_ SUMB_10__5_ NETTRAN_DUMMY_11643 
+ NETTRAN_DUMMY_11644 FA_X1 
XS2_10_4 ab_10__4_ CARRYB_9__4_ SUMB_9__5_ CARRYB_10__4_ SUMB_10__4_ NETTRAN_DUMMY_11645 
+ NETTRAN_DUMMY_11646 FA_X1 
XS2_10_3 ab_10__3_ CARRYB_9__3_ SUMB_9__4_ CARRYB_10__3_ SUMB_10__3_ NETTRAN_DUMMY_11647 
+ NETTRAN_DUMMY_11648 FA_X1 
XS2_10_2 ab_10__2_ CARRYB_9__2_ SUMB_9__3_ CARRYB_10__2_ SUMB_10__2_ NETTRAN_DUMMY_11649 
+ NETTRAN_DUMMY_11650 FA_X1 
XS2_10_1 ab_10__1_ CARRYB_9__1_ SUMB_9__2_ CARRYB_10__1_ SUMB_10__1_ NETTRAN_DUMMY_11651 
+ NETTRAN_DUMMY_11652 FA_X1 
XS1_10_0 ab_10__0_ CARRYB_9__0_ SUMB_9__1_ CARRYB_10__0_ A1_8_ NETTRAN_DUMMY_11653 
+ NETTRAN_DUMMY_11654 FA_X1 
XS3_11_16 ab_11__16_ CARRYB_10__16_ ab_10__17_ CARRYB_11__16_ SUMB_11__16_ NETTRAN_DUMMY_11655 
+ NETTRAN_DUMMY_11656 FA_X1 
XS2_11_15 ab_11__15_ CARRYB_10__15_ SUMB_10__16_ CARRYB_11__15_ SUMB_11__15_ NETTRAN_DUMMY_11657 
+ NETTRAN_DUMMY_11658 FA_X1 
XS2_11_14 ab_11__14_ CARRYB_10__14_ SUMB_10__15_ CARRYB_11__14_ SUMB_11__14_ NETTRAN_DUMMY_11659 
+ NETTRAN_DUMMY_11660 FA_X1 
XS2_11_13 ab_11__13_ CARRYB_10__13_ SUMB_10__14_ CARRYB_11__13_ SUMB_11__13_ NETTRAN_DUMMY_11661 
+ NETTRAN_DUMMY_11662 FA_X1 
XS2_11_12 ab_11__12_ CARRYB_10__12_ SUMB_10__13_ CARRYB_11__12_ SUMB_11__12_ NETTRAN_DUMMY_11663 
+ NETTRAN_DUMMY_11664 FA_X1 
XS2_11_11 ab_11__11_ CARRYB_10__11_ SUMB_10__12_ CARRYB_11__11_ SUMB_11__11_ NETTRAN_DUMMY_11665 
+ NETTRAN_DUMMY_11666 FA_X1 
XS2_11_10 ab_11__10_ CARRYB_10__10_ SUMB_10__11_ CARRYB_11__10_ SUMB_11__10_ NETTRAN_DUMMY_11667 
+ NETTRAN_DUMMY_11668 FA_X1 
XS2_11_9 ab_11__9_ CARRYB_10__9_ SUMB_10__10_ CARRYB_11__9_ SUMB_11__9_ NETTRAN_DUMMY_11669 
+ NETTRAN_DUMMY_11670 FA_X1 
XU26 ab_1__8_ ab_0__9_ n26 NETTRAN_DUMMY_11671 NETTRAN_DUMMY_11672 XOR2_X1 
XU25 ab_1__9_ ab_0__10_ n25 NETTRAN_DUMMY_11673 NETTRAN_DUMMY_11674 XOR2_X1 
XU24 ab_1__10_ ab_0__11_ n24 NETTRAN_DUMMY_11675 NETTRAN_DUMMY_11676 XOR2_X1 
XU23 ab_1__11_ ab_0__12_ n23 NETTRAN_DUMMY_11677 NETTRAN_DUMMY_11678 XOR2_X1 
XU22 ab_1__12_ ab_0__13_ n22 NETTRAN_DUMMY_11679 NETTRAN_DUMMY_11680 XOR2_X1 
XU21 ab_1__13_ ab_0__14_ n21 NETTRAN_DUMMY_11681 NETTRAN_DUMMY_11682 XOR2_X1 
XU20 ab_1__14_ ab_0__15_ n20 NETTRAN_DUMMY_11683 NETTRAN_DUMMY_11684 XOR2_X1 
XU19 ab_1__15_ ab_0__16_ n19 NETTRAN_DUMMY_11685 NETTRAN_DUMMY_11686 XOR2_X1 
XU18 ab_0__17_ ab_1__16_ n18 NETTRAN_DUMMY_11687 NETTRAN_DUMMY_11688 AND2_X1 
XU17 ab_0__1_ ab_1__0_ n17 NETTRAN_DUMMY_11689 NETTRAN_DUMMY_11690 AND2_X1 
XU16 ab_0__2_ ab_1__1_ n16 NETTRAN_DUMMY_11691 NETTRAN_DUMMY_11692 AND2_X1 
XU15 ab_0__3_ ab_1__2_ n15 NETTRAN_DUMMY_11693 NETTRAN_DUMMY_11694 AND2_X1 
XU14 ab_0__4_ ab_1__3_ n14 NETTRAN_DUMMY_11695 NETTRAN_DUMMY_11696 AND2_X1 
XU13 ab_0__5_ ab_1__4_ n13 NETTRAN_DUMMY_11697 NETTRAN_DUMMY_11698 AND2_X1 
XU12 ab_0__6_ ab_1__5_ n12 NETTRAN_DUMMY_11699 NETTRAN_DUMMY_11700 AND2_X1 
XU11 ab_0__7_ ab_1__6_ n11 NETTRAN_DUMMY_11701 NETTRAN_DUMMY_11702 AND2_X1 
XU10 ab_0__8_ ab_1__7_ n10 NETTRAN_DUMMY_11703 NETTRAN_DUMMY_11704 AND2_X1 
XU9 ab_0__9_ ab_1__8_ n9 NETTRAN_DUMMY_11705 NETTRAN_DUMMY_11706 AND2_X1 
XU8 ab_0__10_ ab_1__9_ n8 NETTRAN_DUMMY_11707 NETTRAN_DUMMY_11708 AND2_X1 
XU7 ab_0__11_ ab_1__10_ n7 NETTRAN_DUMMY_11709 NETTRAN_DUMMY_11710 AND2_X1 
XU6 ab_0__12_ ab_1__11_ n6 NETTRAN_DUMMY_11711 NETTRAN_DUMMY_11712 AND2_X1 
XU5 ab_0__13_ ab_1__12_ n5 NETTRAN_DUMMY_11713 NETTRAN_DUMMY_11714 AND2_X1 
XU4 ab_0__14_ ab_1__13_ n4 NETTRAN_DUMMY_11715 NETTRAN_DUMMY_11716 AND2_X1 
XU3 ab_0__15_ ab_1__14_ n3 NETTRAN_DUMMY_11717 NETTRAN_DUMMY_11718 AND2_X1 
XU2 ab_0__16_ ab_1__15_ n2 NETTRAN_DUMMY_11719 NETTRAN_DUMMY_11720 AND2_X1 
XS3_2_16 ab_2__16_ n18 ab_1__17_ CARRYB_2__16_ SUMB_2__16_ NETTRAN_DUMMY_11721 NETTRAN_DUMMY_11722 FA_X1 
XS2_2_15 ab_2__15_ n2 n32 CARRYB_2__15_ SUMB_2__15_ NETTRAN_DUMMY_11723 NETTRAN_DUMMY_11724 FA_X1 
XS2_2_14 ab_2__14_ n3 n19 CARRYB_2__14_ SUMB_2__14_ NETTRAN_DUMMY_11725 NETTRAN_DUMMY_11726 FA_X1 
XS2_2_13 ab_2__13_ n4 n20 CARRYB_2__13_ SUMB_2__13_ NETTRAN_DUMMY_11727 NETTRAN_DUMMY_11728 FA_X1 
XS2_2_12 ab_2__12_ n5 n21 CARRYB_2__12_ SUMB_2__12_ NETTRAN_DUMMY_11729 NETTRAN_DUMMY_11730 FA_X1 
XS2_2_11 ab_2__11_ n6 n22 CARRYB_2__11_ SUMB_2__11_ NETTRAN_DUMMY_11731 NETTRAN_DUMMY_11732 FA_X1 
XS2_2_10 ab_2__10_ n7 n23 CARRYB_2__10_ SUMB_2__10_ NETTRAN_DUMMY_11733 NETTRAN_DUMMY_11734 FA_X1 
XS2_2_9 ab_2__9_ n8 n24 CARRYB_2__9_ SUMB_2__9_ NETTRAN_DUMMY_11735 NETTRAN_DUMMY_11736 FA_X1 
XS2_2_8 ab_2__8_ n9 n25 CARRYB_2__8_ SUMB_2__8_ NETTRAN_DUMMY_11737 NETTRAN_DUMMY_11738 FA_X1 
XS2_2_7 ab_2__7_ n10 n26 CARRYB_2__7_ SUMB_2__7_ NETTRAN_DUMMY_11739 NETTRAN_DUMMY_11740 FA_X1 
XS2_2_6 ab_2__6_ n11 n27 CARRYB_2__6_ SUMB_2__6_ NETTRAN_DUMMY_11741 NETTRAN_DUMMY_11742 FA_X1 
XS2_2_5 ab_2__5_ n12 n28 CARRYB_2__5_ SUMB_2__5_ NETTRAN_DUMMY_11743 NETTRAN_DUMMY_11744 FA_X1 
XS2_2_4 ab_2__4_ n13 n29 CARRYB_2__4_ SUMB_2__4_ NETTRAN_DUMMY_11745 NETTRAN_DUMMY_11746 FA_X1 
XS2_2_3 ab_2__3_ n14 n30 CARRYB_2__3_ SUMB_2__3_ NETTRAN_DUMMY_11747 NETTRAN_DUMMY_11748 FA_X1 
XS2_2_2 ab_2__2_ n15 n31 CARRYB_2__2_ SUMB_2__2_ NETTRAN_DUMMY_11749 NETTRAN_DUMMY_11750 FA_X1 
XS2_2_1 ab_2__1_ n16 n33 CARRYB_2__1_ SUMB_2__1_ NETTRAN_DUMMY_11751 NETTRAN_DUMMY_11752 FA_X1 
XS1_2_0 ab_2__0_ n17 n34 CARRYB_2__0_ A1_0_ NETTRAN_DUMMY_11753 NETTRAN_DUMMY_11754 FA_X1 
XS3_3_16 ab_3__16_ CARRYB_2__16_ ab_2__17_ CARRYB_3__16_ SUMB_3__16_ NETTRAN_DUMMY_11755 
+ NETTRAN_DUMMY_11756 FA_X1 
XS2_3_15 ab_3__15_ CARRYB_2__15_ SUMB_2__16_ CARRYB_3__15_ SUMB_3__15_ NETTRAN_DUMMY_11757 
+ NETTRAN_DUMMY_11758 FA_X1 
XS2_3_14 ab_3__14_ CARRYB_2__14_ SUMB_2__15_ CARRYB_3__14_ SUMB_3__14_ NETTRAN_DUMMY_11759 
+ NETTRAN_DUMMY_11760 FA_X1 
XS2_3_13 ab_3__13_ CARRYB_2__13_ SUMB_2__14_ CARRYB_3__13_ SUMB_3__13_ NETTRAN_DUMMY_11761 
+ NETTRAN_DUMMY_11762 FA_X1 
XS2_3_12 ab_3__12_ CARRYB_2__12_ SUMB_2__13_ CARRYB_3__12_ SUMB_3__12_ NETTRAN_DUMMY_11763 
+ NETTRAN_DUMMY_11764 FA_X1 
XS2_3_11 ab_3__11_ CARRYB_2__11_ SUMB_2__12_ CARRYB_3__11_ SUMB_3__11_ NETTRAN_DUMMY_11765 
+ NETTRAN_DUMMY_11766 FA_X1 
XS2_3_10 ab_3__10_ CARRYB_2__10_ SUMB_2__11_ CARRYB_3__10_ SUMB_3__10_ NETTRAN_DUMMY_11767 
+ NETTRAN_DUMMY_11768 FA_X1 
XS2_3_9 ab_3__9_ CARRYB_2__9_ SUMB_2__10_ CARRYB_3__9_ SUMB_3__9_ NETTRAN_DUMMY_11769 
+ NETTRAN_DUMMY_11770 FA_X1 
XS2_3_8 ab_3__8_ CARRYB_2__8_ SUMB_2__9_ CARRYB_3__8_ SUMB_3__8_ NETTRAN_DUMMY_11771 
+ NETTRAN_DUMMY_11772 FA_X1 
XS2_3_7 ab_3__7_ CARRYB_2__7_ SUMB_2__8_ CARRYB_3__7_ SUMB_3__7_ NETTRAN_DUMMY_11773 
+ NETTRAN_DUMMY_11774 FA_X1 
XS2_3_6 ab_3__6_ CARRYB_2__6_ SUMB_2__7_ CARRYB_3__6_ SUMB_3__6_ NETTRAN_DUMMY_11775 
+ NETTRAN_DUMMY_11776 FA_X1 
XS2_3_5 ab_3__5_ CARRYB_2__5_ SUMB_2__6_ CARRYB_3__5_ SUMB_3__5_ NETTRAN_DUMMY_11777 
+ NETTRAN_DUMMY_11778 FA_X1 
XS2_3_4 ab_3__4_ CARRYB_2__4_ SUMB_2__5_ CARRYB_3__4_ SUMB_3__4_ NETTRAN_DUMMY_11779 
+ NETTRAN_DUMMY_11780 FA_X1 
XS2_3_3 ab_3__3_ CARRYB_2__3_ SUMB_2__4_ CARRYB_3__3_ SUMB_3__3_ NETTRAN_DUMMY_11781 
+ NETTRAN_DUMMY_11782 FA_X1 
XS2_3_2 ab_3__2_ CARRYB_2__2_ SUMB_2__3_ CARRYB_3__2_ SUMB_3__2_ NETTRAN_DUMMY_11783 
+ NETTRAN_DUMMY_11784 FA_X1 
XS2_3_1 ab_3__1_ CARRYB_2__1_ SUMB_2__2_ CARRYB_3__1_ SUMB_3__1_ NETTRAN_DUMMY_11785 
+ NETTRAN_DUMMY_11786 FA_X1 
XS1_3_0 ab_3__0_ CARRYB_2__0_ SUMB_2__1_ CARRYB_3__0_ A1_1_ NETTRAN_DUMMY_11787 
+ NETTRAN_DUMMY_11788 FA_X1 
XS3_4_16 ab_4__16_ CARRYB_3__16_ ab_3__17_ CARRYB_4__16_ SUMB_4__16_ NETTRAN_DUMMY_11789 
+ NETTRAN_DUMMY_11790 FA_X1 
XS2_4_15 ab_4__15_ CARRYB_3__15_ SUMB_3__16_ CARRYB_4__15_ SUMB_4__15_ NETTRAN_DUMMY_11791 
+ NETTRAN_DUMMY_11792 FA_X1 
XS2_4_14 ab_4__14_ CARRYB_3__14_ SUMB_3__15_ CARRYB_4__14_ SUMB_4__14_ NETTRAN_DUMMY_11793 
+ NETTRAN_DUMMY_11794 FA_X1 
XS2_4_13 ab_4__13_ CARRYB_3__13_ SUMB_3__14_ CARRYB_4__13_ SUMB_4__13_ NETTRAN_DUMMY_11795 
+ NETTRAN_DUMMY_11796 FA_X1 
XS2_4_12 ab_4__12_ CARRYB_3__12_ SUMB_3__13_ CARRYB_4__12_ SUMB_4__12_ NETTRAN_DUMMY_11797 
+ NETTRAN_DUMMY_11798 FA_X1 
XS2_4_11 ab_4__11_ CARRYB_3__11_ SUMB_3__12_ CARRYB_4__11_ SUMB_4__11_ NETTRAN_DUMMY_11799 
+ NETTRAN_DUMMY_11800 FA_X1 
XS2_4_10 ab_4__10_ CARRYB_3__10_ SUMB_3__11_ CARRYB_4__10_ SUMB_4__10_ NETTRAN_DUMMY_11801 
+ NETTRAN_DUMMY_11802 FA_X1 
XS2_4_9 ab_4__9_ CARRYB_3__9_ SUMB_3__10_ CARRYB_4__9_ SUMB_4__9_ NETTRAN_DUMMY_11803 
+ NETTRAN_DUMMY_11804 FA_X1 
XS2_4_8 ab_4__8_ CARRYB_3__8_ SUMB_3__9_ CARRYB_4__8_ SUMB_4__8_ NETTRAN_DUMMY_11805 
+ NETTRAN_DUMMY_11806 FA_X1 
XS2_4_7 ab_4__7_ CARRYB_3__7_ SUMB_3__8_ CARRYB_4__7_ SUMB_4__7_ NETTRAN_DUMMY_11807 
+ NETTRAN_DUMMY_11808 FA_X1 
XS2_4_6 ab_4__6_ CARRYB_3__6_ SUMB_3__7_ CARRYB_4__6_ SUMB_4__6_ NETTRAN_DUMMY_11809 
+ NETTRAN_DUMMY_11810 FA_X1 
XS2_4_5 ab_4__5_ CARRYB_3__5_ SUMB_3__6_ CARRYB_4__5_ SUMB_4__5_ NETTRAN_DUMMY_11811 
+ NETTRAN_DUMMY_11812 FA_X1 
XS2_4_4 ab_4__4_ CARRYB_3__4_ SUMB_3__5_ CARRYB_4__4_ SUMB_4__4_ NETTRAN_DUMMY_11813 
+ NETTRAN_DUMMY_11814 FA_X1 
XS2_4_3 ab_4__3_ CARRYB_3__3_ SUMB_3__4_ CARRYB_4__3_ SUMB_4__3_ NETTRAN_DUMMY_11815 
+ NETTRAN_DUMMY_11816 FA_X1 
XS2_4_2 ab_4__2_ CARRYB_3__2_ SUMB_3__3_ CARRYB_4__2_ SUMB_4__2_ NETTRAN_DUMMY_11817 
+ NETTRAN_DUMMY_11818 FA_X1 
XS2_4_1 ab_4__1_ CARRYB_3__1_ SUMB_3__2_ CARRYB_4__1_ SUMB_4__1_ NETTRAN_DUMMY_11819 
+ NETTRAN_DUMMY_11820 FA_X1 
XS1_4_0 ab_4__0_ CARRYB_3__0_ SUMB_3__1_ CARRYB_4__0_ A1_2_ NETTRAN_DUMMY_11821 
+ NETTRAN_DUMMY_11822 FA_X1 
XS3_5_16 ab_5__16_ CARRYB_4__16_ ab_4__17_ CARRYB_5__16_ SUMB_5__16_ NETTRAN_DUMMY_11823 
+ NETTRAN_DUMMY_11824 FA_X1 
XS2_5_15 ab_5__15_ CARRYB_4__15_ SUMB_4__16_ CARRYB_5__15_ SUMB_5__15_ NETTRAN_DUMMY_11825 
+ NETTRAN_DUMMY_11826 FA_X1 
XS2_5_14 ab_5__14_ CARRYB_4__14_ SUMB_4__15_ CARRYB_5__14_ SUMB_5__14_ NETTRAN_DUMMY_11827 
+ NETTRAN_DUMMY_11828 FA_X1 
XS2_5_13 ab_5__13_ CARRYB_4__13_ SUMB_4__14_ CARRYB_5__13_ SUMB_5__13_ NETTRAN_DUMMY_11829 
+ NETTRAN_DUMMY_11830 FA_X1 
XS2_5_12 ab_5__12_ CARRYB_4__12_ SUMB_4__13_ CARRYB_5__12_ SUMB_5__12_ NETTRAN_DUMMY_11831 
+ NETTRAN_DUMMY_11832 FA_X1 
XS2_5_11 ab_5__11_ CARRYB_4__11_ SUMB_4__12_ CARRYB_5__11_ SUMB_5__11_ NETTRAN_DUMMY_11833 
+ NETTRAN_DUMMY_11834 FA_X1 
XS2_5_10 ab_5__10_ CARRYB_4__10_ SUMB_4__11_ CARRYB_5__10_ SUMB_5__10_ NETTRAN_DUMMY_11835 
+ NETTRAN_DUMMY_11836 FA_X1 
XS2_5_9 ab_5__9_ CARRYB_4__9_ SUMB_4__10_ CARRYB_5__9_ SUMB_5__9_ NETTRAN_DUMMY_11837 
+ NETTRAN_DUMMY_11838 FA_X1 
XS2_5_8 ab_5__8_ CARRYB_4__8_ SUMB_4__9_ CARRYB_5__8_ SUMB_5__8_ NETTRAN_DUMMY_11839 
+ NETTRAN_DUMMY_11840 FA_X1 
XS2_5_7 ab_5__7_ CARRYB_4__7_ SUMB_4__8_ CARRYB_5__7_ SUMB_5__7_ NETTRAN_DUMMY_11841 
+ NETTRAN_DUMMY_11842 FA_X1 
XS2_5_6 ab_5__6_ CARRYB_4__6_ SUMB_4__7_ CARRYB_5__6_ SUMB_5__6_ NETTRAN_DUMMY_11843 
+ NETTRAN_DUMMY_11844 FA_X1 
XS2_5_5 ab_5__5_ CARRYB_4__5_ SUMB_4__6_ CARRYB_5__5_ SUMB_5__5_ NETTRAN_DUMMY_11845 
+ NETTRAN_DUMMY_11846 FA_X1 
XS2_5_4 ab_5__4_ CARRYB_4__4_ SUMB_4__5_ CARRYB_5__4_ SUMB_5__4_ NETTRAN_DUMMY_11847 
+ NETTRAN_DUMMY_11848 FA_X1 
XS2_5_3 ab_5__3_ CARRYB_4__3_ SUMB_4__4_ CARRYB_5__3_ SUMB_5__3_ NETTRAN_DUMMY_11849 
+ NETTRAN_DUMMY_11850 FA_X1 
XS2_5_2 ab_5__2_ CARRYB_4__2_ SUMB_4__3_ CARRYB_5__2_ SUMB_5__2_ NETTRAN_DUMMY_11851 
+ NETTRAN_DUMMY_11852 FA_X1 
XS2_5_1 ab_5__1_ CARRYB_4__1_ SUMB_4__2_ CARRYB_5__1_ SUMB_5__1_ NETTRAN_DUMMY_11853 
+ NETTRAN_DUMMY_11854 FA_X1 
XS1_5_0 ab_5__0_ CARRYB_4__0_ SUMB_4__1_ CARRYB_5__0_ A1_3_ NETTRAN_DUMMY_11855 
+ NETTRAN_DUMMY_11856 FA_X1 
XU119 n75 n90 ab_9__12_ NETTRAN_DUMMY_11857 NETTRAN_DUMMY_11858 NOR2_X1 
XU118 n75 n89 ab_9__13_ NETTRAN_DUMMY_11859 NETTRAN_DUMMY_11860 NOR2_X1 
XU117 n75 n88 ab_9__14_ NETTRAN_DUMMY_11861 NETTRAN_DUMMY_11862 NOR2_X1 
XU116 n75 n87 ab_9__15_ NETTRAN_DUMMY_11863 NETTRAN_DUMMY_11864 NOR2_X1 
XU115 n75 n86 ab_9__16_ NETTRAN_DUMMY_11865 NETTRAN_DUMMY_11866 NOR2_X1 
XU114 A[9] n85 ab_9__17_ NETTRAN_DUMMY_11867 NETTRAN_DUMMY_11868 NOR2_X1 
XU113 n75 n101 ab_9__1_ NETTRAN_DUMMY_11869 NETTRAN_DUMMY_11870 NOR2_X1 
XU112 n75 n100 ab_9__2_ NETTRAN_DUMMY_11871 NETTRAN_DUMMY_11872 NOR2_X1 
XU111 n75 n99 ab_9__3_ NETTRAN_DUMMY_11873 NETTRAN_DUMMY_11874 NOR2_X1 
XU110 n75 n98 ab_9__4_ NETTRAN_DUMMY_11875 NETTRAN_DUMMY_11876 NOR2_X1 
XU109 n75 n97 ab_9__5_ NETTRAN_DUMMY_11877 NETTRAN_DUMMY_11878 NOR2_X1 
XU108 n75 n96 ab_9__6_ NETTRAN_DUMMY_11879 NETTRAN_DUMMY_11880 NOR2_X1 
XU107 n75 n95 ab_9__7_ NETTRAN_DUMMY_11881 NETTRAN_DUMMY_11882 NOR2_X1 
XU106 n75 n94 ab_9__8_ NETTRAN_DUMMY_11883 NETTRAN_DUMMY_11884 NOR2_X1 
XU105 n75 n93 ab_9__9_ NETTRAN_DUMMY_11885 NETTRAN_DUMMY_11886 NOR2_X1 
XU103 B[0] n102 NETTRAN_DUMMY_11887 NETTRAN_DUMMY_11888 INV_X1 
XU102 B[1] n101 NETTRAN_DUMMY_11889 NETTRAN_DUMMY_11890 INV_X1 
XU101 A[15] SUMB_15__0_ n69 NETTRAN_DUMMY_11891 NETTRAN_DUMMY_11892 XOR2_X1 
XU100 B[2] n100 NETTRAN_DUMMY_11893 NETTRAN_DUMMY_11894 INV_X1 
XU99 B[3] n99 NETTRAN_DUMMY_11895 NETTRAN_DUMMY_11896 INV_X1 
XU98 B[4] n98 NETTRAN_DUMMY_11897 NETTRAN_DUMMY_11898 INV_X1 
XU97 B[5] n97 NETTRAN_DUMMY_11899 NETTRAN_DUMMY_11900 INV_X1 
XU96 B[6] n96 NETTRAN_DUMMY_11901 NETTRAN_DUMMY_11902 INV_X1 
XU95 B[7] n95 NETTRAN_DUMMY_11903 NETTRAN_DUMMY_11904 INV_X1 
XU94 B[8] n94 NETTRAN_DUMMY_11905 NETTRAN_DUMMY_11906 INV_X1 
XU93 B[9] n93 NETTRAN_DUMMY_11907 NETTRAN_DUMMY_11908 INV_X1 
XU92 B[10] n92 NETTRAN_DUMMY_11909 NETTRAN_DUMMY_11910 INV_X1 
XU91 B[11] n91 NETTRAN_DUMMY_11911 NETTRAN_DUMMY_11912 INV_X1 
XU90 B[12] n90 NETTRAN_DUMMY_11913 NETTRAN_DUMMY_11914 INV_X1 
XU89 A[15] SUMB_15__0_ n68 NETTRAN_DUMMY_11915 NETTRAN_DUMMY_11916 AND2_X1 
XU88 B[13] n89 NETTRAN_DUMMY_11917 NETTRAN_DUMMY_11918 INV_X1 
XU87 B[14] n88 NETTRAN_DUMMY_11919 NETTRAN_DUMMY_11920 INV_X1 
XU86 B[15] n87 NETTRAN_DUMMY_11921 NETTRAN_DUMMY_11922 INV_X1 
XU85 B[16] n86 NETTRAN_DUMMY_11923 NETTRAN_DUMMY_11924 INV_X1 
XU84 B[17] n85 NETTRAN_DUMMY_11925 NETTRAN_DUMMY_11926 INV_X1 
XU83 A[0] n84 NETTRAN_DUMMY_11927 NETTRAN_DUMMY_11928 INV_X1 
XU82 A[1] n83 NETTRAN_DUMMY_11929 NETTRAN_DUMMY_11930 INV_X1 
XU81 A[2] n82 NETTRAN_DUMMY_11931 NETTRAN_DUMMY_11932 INV_X1 
XU80 A[3] n81 NETTRAN_DUMMY_11933 NETTRAN_DUMMY_11934 INV_X1 
XU79 A[4] n80 NETTRAN_DUMMY_11935 NETTRAN_DUMMY_11936 INV_X1 
XU78 A[5] n79 NETTRAN_DUMMY_11937 NETTRAN_DUMMY_11938 INV_X1 
XU77 A[6] n78 NETTRAN_DUMMY_11939 NETTRAN_DUMMY_11940 INV_X1 
XU76 A[7] n77 NETTRAN_DUMMY_11941 NETTRAN_DUMMY_11942 INV_X1 
XU75 A[8] n76 NETTRAN_DUMMY_11943 NETTRAN_DUMMY_11944 INV_X1 
XU74 A[9] n75 NETTRAN_DUMMY_11945 NETTRAN_DUMMY_11946 INV_X1 
XU73 A[10] n74 NETTRAN_DUMMY_11947 NETTRAN_DUMMY_11948 INV_X1 
XU72 A[11] n73 NETTRAN_DUMMY_11949 NETTRAN_DUMMY_11950 INV_X1 
XU71 A[12] n72 NETTRAN_DUMMY_11951 NETTRAN_DUMMY_11952 INV_X1 
XU70 A[13] n71 NETTRAN_DUMMY_11953 NETTRAN_DUMMY_11954 INV_X1 
XU69 A[14] n35 NETTRAN_DUMMY_11955 NETTRAN_DUMMY_11956 INV_X1 
XU68 CARRYB_15__15_ SUMB_15__16_ n67 NETTRAN_DUMMY_11957 NETTRAN_DUMMY_11958 XOR2_X1 
XU67 CARRYB_15__13_ SUMB_15__14_ n66 NETTRAN_DUMMY_11959 NETTRAN_DUMMY_11960 XOR2_X1 
XU66 CARRYB_15__11_ SUMB_15__12_ n65 NETTRAN_DUMMY_11961 NETTRAN_DUMMY_11962 XOR2_X1 
XU65 CARRYB_15__9_ SUMB_15__10_ n64 NETTRAN_DUMMY_11963 NETTRAN_DUMMY_11964 XOR2_X1 
XU64 CARRYB_15__7_ SUMB_15__8_ n63 NETTRAN_DUMMY_11965 NETTRAN_DUMMY_11966 XOR2_X1 
XU63 CARRYB_15__5_ SUMB_15__6_ n62 NETTRAN_DUMMY_11967 NETTRAN_DUMMY_11968 XOR2_X1 
XU62 CARRYB_15__15_ SUMB_15__16_ n61 NETTRAN_DUMMY_11969 NETTRAN_DUMMY_11970 AND2_X1 
XU61 CARRYB_15__14_ SUMB_15__15_ n60 NETTRAN_DUMMY_11971 NETTRAN_DUMMY_11972 AND2_X1 
XU60 CARRYB_15__13_ SUMB_15__14_ n59 NETTRAN_DUMMY_11973 NETTRAN_DUMMY_11974 AND2_X1 
XU59 CARRYB_15__12_ SUMB_15__13_ n58 NETTRAN_DUMMY_11975 NETTRAN_DUMMY_11976 AND2_X1 
XU58 CARRYB_15__11_ SUMB_15__12_ n57 NETTRAN_DUMMY_11977 NETTRAN_DUMMY_11978 AND2_X1 
XU57 CARRYB_15__10_ SUMB_15__11_ n56 NETTRAN_DUMMY_11979 NETTRAN_DUMMY_11980 AND2_X1 
XU56 CARRYB_15__9_ SUMB_15__10_ n55 NETTRAN_DUMMY_11981 NETTRAN_DUMMY_11982 AND2_X1 
XU55 CARRYB_15__8_ SUMB_15__9_ n54 NETTRAN_DUMMY_11983 NETTRAN_DUMMY_11984 AND2_X1 
XU54 CARRYB_15__7_ SUMB_15__8_ n53 NETTRAN_DUMMY_11985 NETTRAN_DUMMY_11986 AND2_X1 
XU53 CARRYB_15__6_ SUMB_15__7_ n52 NETTRAN_DUMMY_11987 NETTRAN_DUMMY_11988 AND2_X1 
XU52 CARRYB_15__5_ SUMB_15__6_ n51 NETTRAN_DUMMY_11989 NETTRAN_DUMMY_11990 AND2_X1 
XU51 CARRYB_15__4_ SUMB_15__5_ n50 NETTRAN_DUMMY_11991 NETTRAN_DUMMY_11992 AND2_X1 
XU50 CARRYB_15__16_ SUMB_15__17_ n49 NETTRAN_DUMMY_11993 NETTRAN_DUMMY_11994 AND2_X1 
XU49 CARRYB_15__16_ SUMB_15__17_ n48 NETTRAN_DUMMY_11995 NETTRAN_DUMMY_11996 XOR2_X1 
XU48 CARRYB_15__14_ SUMB_15__15_ n47 NETTRAN_DUMMY_11997 NETTRAN_DUMMY_11998 XOR2_X1 
XU47 CARRYB_15__12_ SUMB_15__13_ n46 NETTRAN_DUMMY_11999 NETTRAN_DUMMY_12000 XOR2_X1 
XU46 CARRYB_15__10_ SUMB_15__11_ n45 NETTRAN_DUMMY_12001 NETTRAN_DUMMY_12002 XOR2_X1 
XU45 CARRYB_15__8_ SUMB_15__9_ n44 NETTRAN_DUMMY_12003 NETTRAN_DUMMY_12004 XOR2_X1 
XU44 CARRYB_15__6_ SUMB_15__7_ n43 NETTRAN_DUMMY_12005 NETTRAN_DUMMY_12006 XOR2_X1 
XU43 CARRYB_15__3_ SUMB_15__4_ n42 NETTRAN_DUMMY_12007 NETTRAN_DUMMY_12008 XOR2_X1 
XU42 CARRYB_15__3_ SUMB_15__4_ n41 NETTRAN_DUMMY_12009 NETTRAN_DUMMY_12010 AND2_X1 
XU41 CARRYB_15__2_ SUMB_15__3_ n40 NETTRAN_DUMMY_12011 NETTRAN_DUMMY_12012 AND2_X1 
XU40 CARRYB_15__0_ SUMB_15__1_ n39 NETTRAN_DUMMY_12013 NETTRAN_DUMMY_12014 AND2_X1 
XU39 CARRYB_15__0_ SUMB_15__1_ n38 NETTRAN_DUMMY_12015 NETTRAN_DUMMY_12016 XOR2_X1 
XU38 CARRYB_15__4_ SUMB_15__5_ n37 NETTRAN_DUMMY_12017 NETTRAN_DUMMY_12018 XOR2_X1 
XU37 CARRYB_15__2_ SUMB_15__3_ n36 NETTRAN_DUMMY_12019 NETTRAN_DUMMY_12020 XOR2_X1 
XU36 ab_1__0_ ab_0__1_ n158 NETTRAN_DUMMY_12021 NETTRAN_DUMMY_12022 XOR2_X1 
XU35 CARRYB_15__17_ n70 NETTRAN_DUMMY_12023 NETTRAN_DUMMY_12024 INV_X1 
XU34 ab_1__1_ ab_0__2_ n34 NETTRAN_DUMMY_12025 NETTRAN_DUMMY_12026 XOR2_X1 
XU33 ab_1__2_ ab_0__3_ n33 NETTRAN_DUMMY_12027 NETTRAN_DUMMY_12028 XOR2_X1 
XU32 ab_1__16_ ab_0__17_ n32 NETTRAN_DUMMY_12029 NETTRAN_DUMMY_12030 XOR2_X1 
XU31 ab_1__3_ ab_0__4_ n31 NETTRAN_DUMMY_12031 NETTRAN_DUMMY_12032 XOR2_X1 
XU30 ab_1__4_ ab_0__5_ n30 NETTRAN_DUMMY_12033 NETTRAN_DUMMY_12034 XOR2_X1 
XU29 ab_1__5_ ab_0__6_ n29 NETTRAN_DUMMY_12035 NETTRAN_DUMMY_12036 XOR2_X1 
XU28 ab_1__6_ ab_0__7_ n28 NETTRAN_DUMMY_12037 NETTRAN_DUMMY_12038 XOR2_X1 
XU27 ab_1__7_ ab_0__8_ n27 NETTRAN_DUMMY_12039 NETTRAN_DUMMY_12040 XOR2_X1 
XU212 n156 n80 ab_4__0_ NETTRAN_DUMMY_12041 NETTRAN_DUMMY_12042 NOR2_X1 
XU211 n92 n80 ab_4__10_ NETTRAN_DUMMY_12043 NETTRAN_DUMMY_12044 NOR2_X1 
XU210 n91 n80 ab_4__11_ NETTRAN_DUMMY_12045 NETTRAN_DUMMY_12046 NOR2_X1 
XU209 n90 n80 ab_4__12_ NETTRAN_DUMMY_12047 NETTRAN_DUMMY_12048 NOR2_X1 
XU208 n89 n80 ab_4__13_ NETTRAN_DUMMY_12049 NETTRAN_DUMMY_12050 NOR2_X1 
XU207 n88 n80 ab_4__14_ NETTRAN_DUMMY_12051 NETTRAN_DUMMY_12052 NOR2_X1 
XU206 n87 n80 ab_4__15_ NETTRAN_DUMMY_12053 NETTRAN_DUMMY_12054 NOR2_X1 
XU205 n86 n80 ab_4__16_ NETTRAN_DUMMY_12055 NETTRAN_DUMMY_12056 NOR2_X1 
XU204 A[4] n85 ab_4__17_ NETTRAN_DUMMY_12057 NETTRAN_DUMMY_12058 NOR2_X1 
XU203 n101 n80 ab_4__1_ NETTRAN_DUMMY_12059 NETTRAN_DUMMY_12060 NOR2_X1 
XU202 n100 n80 ab_4__2_ NETTRAN_DUMMY_12061 NETTRAN_DUMMY_12062 NOR2_X1 
XU201 n99 n80 ab_4__3_ NETTRAN_DUMMY_12063 NETTRAN_DUMMY_12064 NOR2_X1 
XU200 n98 n80 ab_4__4_ NETTRAN_DUMMY_12065 NETTRAN_DUMMY_12066 NOR2_X1 
XU199 n97 n80 ab_4__5_ NETTRAN_DUMMY_12067 NETTRAN_DUMMY_12068 NOR2_X1 
XU198 n96 n80 ab_4__6_ NETTRAN_DUMMY_12069 NETTRAN_DUMMY_12070 NOR2_X1 
XU197 n95 n80 ab_4__7_ NETTRAN_DUMMY_12071 NETTRAN_DUMMY_12072 NOR2_X1 
XU196 n94 n80 ab_4__8_ NETTRAN_DUMMY_12073 NETTRAN_DUMMY_12074 NOR2_X1 
XU195 n93 n80 ab_4__9_ NETTRAN_DUMMY_12075 NETTRAN_DUMMY_12076 NOR2_X1 
XU194 n156 n79 ab_5__0_ NETTRAN_DUMMY_12077 NETTRAN_DUMMY_12078 NOR2_X1 
XU193 n92 n79 ab_5__10_ NETTRAN_DUMMY_12079 NETTRAN_DUMMY_12080 NOR2_X1 
XU192 n91 n79 ab_5__11_ NETTRAN_DUMMY_12081 NETTRAN_DUMMY_12082 NOR2_X1 
XU191 n90 n79 ab_5__12_ NETTRAN_DUMMY_12083 NETTRAN_DUMMY_12084 NOR2_X1 
XU190 n89 n79 ab_5__13_ NETTRAN_DUMMY_12085 NETTRAN_DUMMY_12086 NOR2_X1 
XU189 n88 n79 ab_5__14_ NETTRAN_DUMMY_12087 NETTRAN_DUMMY_12088 NOR2_X1 
XU188 n87 n79 ab_5__15_ NETTRAN_DUMMY_12089 NETTRAN_DUMMY_12090 NOR2_X1 
XU187 n86 n79 ab_5__16_ NETTRAN_DUMMY_12091 NETTRAN_DUMMY_12092 NOR2_X1 
XU186 A[5] n85 ab_5__17_ NETTRAN_DUMMY_12093 NETTRAN_DUMMY_12094 NOR2_X1 
XU185 n101 n79 ab_5__1_ NETTRAN_DUMMY_12095 NETTRAN_DUMMY_12096 NOR2_X1 
XU184 n100 n79 ab_5__2_ NETTRAN_DUMMY_12097 NETTRAN_DUMMY_12098 NOR2_X1 
XU183 n99 n79 ab_5__3_ NETTRAN_DUMMY_12099 NETTRAN_DUMMY_12100 NOR2_X1 
XU182 n98 n79 ab_5__4_ NETTRAN_DUMMY_12101 NETTRAN_DUMMY_12102 NOR2_X1 
XU181 n97 n79 ab_5__5_ NETTRAN_DUMMY_12103 NETTRAN_DUMMY_12104 NOR2_X1 
XU180 n96 n79 ab_5__6_ NETTRAN_DUMMY_12105 NETTRAN_DUMMY_12106 NOR2_X1 
XU179 n95 n79 ab_5__7_ NETTRAN_DUMMY_12107 NETTRAN_DUMMY_12108 NOR2_X1 
XU178 n94 n79 ab_5__8_ NETTRAN_DUMMY_12109 NETTRAN_DUMMY_12110 NOR2_X1 
XU177 n93 n79 ab_5__9_ NETTRAN_DUMMY_12111 NETTRAN_DUMMY_12112 NOR2_X1 
XU176 n156 n78 ab_6__0_ NETTRAN_DUMMY_12113 NETTRAN_DUMMY_12114 NOR2_X1 
XU175 n92 n78 ab_6__10_ NETTRAN_DUMMY_12115 NETTRAN_DUMMY_12116 NOR2_X1 
XU174 n91 n78 ab_6__11_ NETTRAN_DUMMY_12117 NETTRAN_DUMMY_12118 NOR2_X1 
XU173 n90 n78 ab_6__12_ NETTRAN_DUMMY_12119 NETTRAN_DUMMY_12120 NOR2_X1 
XU172 n89 n78 ab_6__13_ NETTRAN_DUMMY_12121 NETTRAN_DUMMY_12122 NOR2_X1 
XU171 n88 n78 ab_6__14_ NETTRAN_DUMMY_12123 NETTRAN_DUMMY_12124 NOR2_X1 
XU170 n87 n78 ab_6__15_ NETTRAN_DUMMY_12125 NETTRAN_DUMMY_12126 NOR2_X1 
XU169 n86 n78 ab_6__16_ NETTRAN_DUMMY_12127 NETTRAN_DUMMY_12128 NOR2_X1 
XU168 A[6] n85 ab_6__17_ NETTRAN_DUMMY_12129 NETTRAN_DUMMY_12130 NOR2_X1 
XU167 n101 n78 ab_6__1_ NETTRAN_DUMMY_12131 NETTRAN_DUMMY_12132 NOR2_X1 
XU166 n100 n78 ab_6__2_ NETTRAN_DUMMY_12133 NETTRAN_DUMMY_12134 NOR2_X1 
XU165 n99 n78 ab_6__3_ NETTRAN_DUMMY_12135 NETTRAN_DUMMY_12136 NOR2_X1 
XU164 n98 n78 ab_6__4_ NETTRAN_DUMMY_12137 NETTRAN_DUMMY_12138 NOR2_X1 
XU163 n97 n78 ab_6__5_ NETTRAN_DUMMY_12139 NETTRAN_DUMMY_12140 NOR2_X1 
XU162 n96 n78 ab_6__6_ NETTRAN_DUMMY_12141 NETTRAN_DUMMY_12142 NOR2_X1 
XU161 n95 n78 ab_6__7_ NETTRAN_DUMMY_12143 NETTRAN_DUMMY_12144 NOR2_X1 
XU160 n94 n78 ab_6__8_ NETTRAN_DUMMY_12145 NETTRAN_DUMMY_12146 NOR2_X1 
XU159 n93 n78 ab_6__9_ NETTRAN_DUMMY_12147 NETTRAN_DUMMY_12148 NOR2_X1 
XU158 n156 n77 ab_7__0_ NETTRAN_DUMMY_12149 NETTRAN_DUMMY_12150 NOR2_X1 
XU157 n92 n77 ab_7__10_ NETTRAN_DUMMY_12151 NETTRAN_DUMMY_12152 NOR2_X1 
XU156 n91 n77 ab_7__11_ NETTRAN_DUMMY_12153 NETTRAN_DUMMY_12154 NOR2_X1 
XU155 n90 n77 ab_7__12_ NETTRAN_DUMMY_12155 NETTRAN_DUMMY_12156 NOR2_X1 
XU154 n89 n77 ab_7__13_ NETTRAN_DUMMY_12157 NETTRAN_DUMMY_12158 NOR2_X1 
XU153 n88 n77 ab_7__14_ NETTRAN_DUMMY_12159 NETTRAN_DUMMY_12160 NOR2_X1 
XU152 n87 n77 ab_7__15_ NETTRAN_DUMMY_12161 NETTRAN_DUMMY_12162 NOR2_X1 
XU151 n86 n77 ab_7__16_ NETTRAN_DUMMY_12163 NETTRAN_DUMMY_12164 NOR2_X1 
XU150 A[7] n85 ab_7__17_ NETTRAN_DUMMY_12165 NETTRAN_DUMMY_12166 NOR2_X1 
XU149 n101 n77 ab_7__1_ NETTRAN_DUMMY_12167 NETTRAN_DUMMY_12168 NOR2_X1 
XU148 n100 n77 ab_7__2_ NETTRAN_DUMMY_12169 NETTRAN_DUMMY_12170 NOR2_X1 
XU147 n99 n77 ab_7__3_ NETTRAN_DUMMY_12171 NETTRAN_DUMMY_12172 NOR2_X1 
XU146 n98 n77 ab_7__4_ NETTRAN_DUMMY_12173 NETTRAN_DUMMY_12174 NOR2_X1 
XU145 n97 n77 ab_7__5_ NETTRAN_DUMMY_12175 NETTRAN_DUMMY_12176 NOR2_X1 
XU144 n96 n77 ab_7__6_ NETTRAN_DUMMY_12177 NETTRAN_DUMMY_12178 NOR2_X1 
XU143 n95 n77 ab_7__7_ NETTRAN_DUMMY_12179 NETTRAN_DUMMY_12180 NOR2_X1 
XU142 n94 n77 ab_7__8_ NETTRAN_DUMMY_12181 NETTRAN_DUMMY_12182 NOR2_X1 
XU141 n93 n77 ab_7__9_ NETTRAN_DUMMY_12183 NETTRAN_DUMMY_12184 NOR2_X1 
XU140 n156 n76 ab_8__0_ NETTRAN_DUMMY_12185 NETTRAN_DUMMY_12186 NOR2_X1 
XU139 n92 n76 ab_8__10_ NETTRAN_DUMMY_12187 NETTRAN_DUMMY_12188 NOR2_X1 
XU138 n91 n76 ab_8__11_ NETTRAN_DUMMY_12189 NETTRAN_DUMMY_12190 NOR2_X1 
XU137 n90 n76 ab_8__12_ NETTRAN_DUMMY_12191 NETTRAN_DUMMY_12192 NOR2_X1 
XU136 n89 n76 ab_8__13_ NETTRAN_DUMMY_12193 NETTRAN_DUMMY_12194 NOR2_X1 
XU135 n88 n76 ab_8__14_ NETTRAN_DUMMY_12195 NETTRAN_DUMMY_12196 NOR2_X1 
XU134 n87 n76 ab_8__15_ NETTRAN_DUMMY_12197 NETTRAN_DUMMY_12198 NOR2_X1 
XU133 n86 n76 ab_8__16_ NETTRAN_DUMMY_12199 NETTRAN_DUMMY_12200 NOR2_X1 
XU132 A[8] n85 ab_8__17_ NETTRAN_DUMMY_12201 NETTRAN_DUMMY_12202 NOR2_X1 
XU131 n101 n76 ab_8__1_ NETTRAN_DUMMY_12203 NETTRAN_DUMMY_12204 NOR2_X1 
XU130 n100 n76 ab_8__2_ NETTRAN_DUMMY_12205 NETTRAN_DUMMY_12206 NOR2_X1 
XU129 n99 n76 ab_8__3_ NETTRAN_DUMMY_12207 NETTRAN_DUMMY_12208 NOR2_X1 
XU128 n98 n76 ab_8__4_ NETTRAN_DUMMY_12209 NETTRAN_DUMMY_12210 NOR2_X1 
XU127 n97 n76 ab_8__5_ NETTRAN_DUMMY_12211 NETTRAN_DUMMY_12212 NOR2_X1 
XU126 n96 n76 ab_8__6_ NETTRAN_DUMMY_12213 NETTRAN_DUMMY_12214 NOR2_X1 
XU125 n95 n76 ab_8__7_ NETTRAN_DUMMY_12215 NETTRAN_DUMMY_12216 NOR2_X1 
XU124 n94 n76 ab_8__8_ NETTRAN_DUMMY_12217 NETTRAN_DUMMY_12218 NOR2_X1 
XU123 n93 n76 ab_8__9_ NETTRAN_DUMMY_12219 NETTRAN_DUMMY_12220 NOR2_X1 
XU122 n75 n156 ab_9__0_ NETTRAN_DUMMY_12221 NETTRAN_DUMMY_12222 NOR2_X1 
XU121 n75 n92 ab_9__10_ NETTRAN_DUMMY_12223 NETTRAN_DUMMY_12224 NOR2_X1 
XU120 n75 n91 ab_9__11_ NETTRAN_DUMMY_12225 NETTRAN_DUMMY_12226 NOR2_X1 
XU305 n95 n71 ab_13__7_ NETTRAN_DUMMY_12227 NETTRAN_DUMMY_12228 NOR2_X1 
XU304 n94 n71 ab_13__8_ NETTRAN_DUMMY_12229 NETTRAN_DUMMY_12230 NOR2_X1 
XU303 n93 n71 ab_13__9_ NETTRAN_DUMMY_12231 NETTRAN_DUMMY_12232 NOR2_X1 
XU302 n156 n35 ab_14__0_ NETTRAN_DUMMY_12233 NETTRAN_DUMMY_12234 NOR2_X1 
XU301 n92 n35 ab_14__10_ NETTRAN_DUMMY_12235 NETTRAN_DUMMY_12236 NOR2_X1 
XU300 n91 n35 ab_14__11_ NETTRAN_DUMMY_12237 NETTRAN_DUMMY_12238 NOR2_X1 
XU299 n90 n35 ab_14__12_ NETTRAN_DUMMY_12239 NETTRAN_DUMMY_12240 NOR2_X1 
XU298 n89 n35 ab_14__13_ NETTRAN_DUMMY_12241 NETTRAN_DUMMY_12242 NOR2_X1 
XU297 n88 n35 ab_14__14_ NETTRAN_DUMMY_12243 NETTRAN_DUMMY_12244 NOR2_X1 
XU296 n87 n35 ab_14__15_ NETTRAN_DUMMY_12245 NETTRAN_DUMMY_12246 NOR2_X1 
XU295 n86 n35 ab_14__16_ NETTRAN_DUMMY_12247 NETTRAN_DUMMY_12248 NOR2_X1 
XU294 A[14] n85 ab_14__17_ NETTRAN_DUMMY_12249 NETTRAN_DUMMY_12250 NOR2_X1 
XU293 n101 n35 ab_14__1_ NETTRAN_DUMMY_12251 NETTRAN_DUMMY_12252 NOR2_X1 
XU292 n100 n35 ab_14__2_ NETTRAN_DUMMY_12253 NETTRAN_DUMMY_12254 NOR2_X1 
XU291 n99 n35 ab_14__3_ NETTRAN_DUMMY_12255 NETTRAN_DUMMY_12256 NOR2_X1 
XU290 n98 n35 ab_14__4_ NETTRAN_DUMMY_12257 NETTRAN_DUMMY_12258 NOR2_X1 
XU289 n97 n35 ab_14__5_ NETTRAN_DUMMY_12259 NETTRAN_DUMMY_12260 NOR2_X1 
XU288 n96 n35 ab_14__6_ NETTRAN_DUMMY_12261 NETTRAN_DUMMY_12262 NOR2_X1 
XU287 n95 n35 ab_14__7_ NETTRAN_DUMMY_12263 NETTRAN_DUMMY_12264 NOR2_X1 
XU286 n94 n35 ab_14__8_ NETTRAN_DUMMY_12265 NETTRAN_DUMMY_12266 NOR2_X1 
XU285 n93 n35 ab_14__9_ NETTRAN_DUMMY_12267 NETTRAN_DUMMY_12268 NOR2_X1 
XU284 B[0] n1 ab_15__0_ NETTRAN_DUMMY_12269 NETTRAN_DUMMY_12270 NOR2_X1 
XU283 B[10] n1 ab_15__10_ NETTRAN_DUMMY_12271 NETTRAN_DUMMY_12272 NOR2_X1 
XU282 B[11] n1 ab_15__11_ NETTRAN_DUMMY_12273 NETTRAN_DUMMY_12274 NOR2_X1 
XU281 B[12] n1 ab_15__12_ NETTRAN_DUMMY_12275 NETTRAN_DUMMY_12276 NOR2_X1 
XU280 B[13] n1 ab_15__13_ NETTRAN_DUMMY_12277 NETTRAN_DUMMY_12278 NOR2_X1 
XU279 B[14] n1 ab_15__14_ NETTRAN_DUMMY_12279 NETTRAN_DUMMY_12280 NOR2_X1 
XU278 B[15] n1 ab_15__15_ NETTRAN_DUMMY_12281 NETTRAN_DUMMY_12282 NOR2_X1 
XU277 B[16] n1 ab_15__16_ NETTRAN_DUMMY_12283 NETTRAN_DUMMY_12284 NOR2_X1 
XU276 n85 n1 ab_15__17_ NETTRAN_DUMMY_12285 NETTRAN_DUMMY_12286 NOR2_X1 
XU275 B[1] n1 ab_15__1_ NETTRAN_DUMMY_12287 NETTRAN_DUMMY_12288 NOR2_X1 
XU274 B[2] n1 ab_15__2_ NETTRAN_DUMMY_12289 NETTRAN_DUMMY_12290 NOR2_X1 
XU273 B[3] n1 ab_15__3_ NETTRAN_DUMMY_12291 NETTRAN_DUMMY_12292 NOR2_X1 
XU272 B[4] n1 ab_15__4_ NETTRAN_DUMMY_12293 NETTRAN_DUMMY_12294 NOR2_X1 
XU271 B[5] n1 ab_15__5_ NETTRAN_DUMMY_12295 NETTRAN_DUMMY_12296 NOR2_X1 
XU270 B[6] n1 ab_15__6_ NETTRAN_DUMMY_12297 NETTRAN_DUMMY_12298 NOR2_X1 
XU269 B[7] n1 ab_15__7_ NETTRAN_DUMMY_12299 NETTRAN_DUMMY_12300 NOR2_X1 
XU268 B[8] n1 ab_15__8_ NETTRAN_DUMMY_12301 NETTRAN_DUMMY_12302 NOR2_X1 
XU267 B[9] n1 ab_15__9_ NETTRAN_DUMMY_12303 NETTRAN_DUMMY_12304 NOR2_X1 
XU266 n156 n83 ab_1__0_ NETTRAN_DUMMY_12305 NETTRAN_DUMMY_12306 NOR2_X1 
XU265 n92 n83 ab_1__10_ NETTRAN_DUMMY_12307 NETTRAN_DUMMY_12308 NOR2_X1 
XU264 n91 n83 ab_1__11_ NETTRAN_DUMMY_12309 NETTRAN_DUMMY_12310 NOR2_X1 
XU263 n90 n83 ab_1__12_ NETTRAN_DUMMY_12311 NETTRAN_DUMMY_12312 NOR2_X1 
XU262 n89 n83 ab_1__13_ NETTRAN_DUMMY_12313 NETTRAN_DUMMY_12314 NOR2_X1 
XU261 n88 n83 ab_1__14_ NETTRAN_DUMMY_12315 NETTRAN_DUMMY_12316 NOR2_X1 
XU260 n87 n83 ab_1__15_ NETTRAN_DUMMY_12317 NETTRAN_DUMMY_12318 NOR2_X1 
XU259 n86 n83 ab_1__16_ NETTRAN_DUMMY_12319 NETTRAN_DUMMY_12320 NOR2_X1 
XU258 A[1] n85 ab_1__17_ NETTRAN_DUMMY_12321 NETTRAN_DUMMY_12322 NOR2_X1 
XU257 n101 n83 ab_1__1_ NETTRAN_DUMMY_12323 NETTRAN_DUMMY_12324 NOR2_X1 
XU256 n100 n83 ab_1__2_ NETTRAN_DUMMY_12325 NETTRAN_DUMMY_12326 NOR2_X1 
XU255 n99 n83 ab_1__3_ NETTRAN_DUMMY_12327 NETTRAN_DUMMY_12328 NOR2_X1 
XU254 n98 n83 ab_1__4_ NETTRAN_DUMMY_12329 NETTRAN_DUMMY_12330 NOR2_X1 
XU253 n97 n83 ab_1__5_ NETTRAN_DUMMY_12331 NETTRAN_DUMMY_12332 NOR2_X1 
XU252 n96 n83 ab_1__6_ NETTRAN_DUMMY_12333 NETTRAN_DUMMY_12334 NOR2_X1 
XU251 n95 n83 ab_1__7_ NETTRAN_DUMMY_12335 NETTRAN_DUMMY_12336 NOR2_X1 
XU250 n94 n83 ab_1__8_ NETTRAN_DUMMY_12337 NETTRAN_DUMMY_12338 NOR2_X1 
XU249 n93 n83 ab_1__9_ NETTRAN_DUMMY_12339 NETTRAN_DUMMY_12340 NOR2_X1 
XU248 n156 n82 ab_2__0_ NETTRAN_DUMMY_12341 NETTRAN_DUMMY_12342 NOR2_X1 
XU247 n92 n82 ab_2__10_ NETTRAN_DUMMY_12343 NETTRAN_DUMMY_12344 NOR2_X1 
XU246 n91 n82 ab_2__11_ NETTRAN_DUMMY_12345 NETTRAN_DUMMY_12346 NOR2_X1 
XU245 n90 n82 ab_2__12_ NETTRAN_DUMMY_12347 NETTRAN_DUMMY_12348 NOR2_X1 
XU244 n89 n82 ab_2__13_ NETTRAN_DUMMY_12349 NETTRAN_DUMMY_12350 NOR2_X1 
XU243 n88 n82 ab_2__14_ NETTRAN_DUMMY_12351 NETTRAN_DUMMY_12352 NOR2_X1 
XU242 n87 n82 ab_2__15_ NETTRAN_DUMMY_12353 NETTRAN_DUMMY_12354 NOR2_X1 
XU241 n86 n82 ab_2__16_ NETTRAN_DUMMY_12355 NETTRAN_DUMMY_12356 NOR2_X1 
XU240 A[2] n85 ab_2__17_ NETTRAN_DUMMY_12357 NETTRAN_DUMMY_12358 NOR2_X1 
XU239 n101 n82 ab_2__1_ NETTRAN_DUMMY_12359 NETTRAN_DUMMY_12360 NOR2_X1 
XU238 n100 n82 ab_2__2_ NETTRAN_DUMMY_12361 NETTRAN_DUMMY_12362 NOR2_X1 
XU237 n99 n82 ab_2__3_ NETTRAN_DUMMY_12363 NETTRAN_DUMMY_12364 NOR2_X1 
XU236 n98 n82 ab_2__4_ NETTRAN_DUMMY_12365 NETTRAN_DUMMY_12366 NOR2_X1 
XU235 n97 n82 ab_2__5_ NETTRAN_DUMMY_12367 NETTRAN_DUMMY_12368 NOR2_X1 
XU234 n96 n82 ab_2__6_ NETTRAN_DUMMY_12369 NETTRAN_DUMMY_12370 NOR2_X1 
XU233 n95 n82 ab_2__7_ NETTRAN_DUMMY_12371 NETTRAN_DUMMY_12372 NOR2_X1 
XU232 n94 n82 ab_2__8_ NETTRAN_DUMMY_12373 NETTRAN_DUMMY_12374 NOR2_X1 
XU231 n93 n82 ab_2__9_ NETTRAN_DUMMY_12375 NETTRAN_DUMMY_12376 NOR2_X1 
XU230 n156 n81 ab_3__0_ NETTRAN_DUMMY_12377 NETTRAN_DUMMY_12378 NOR2_X1 
XU229 n92 n81 ab_3__10_ NETTRAN_DUMMY_12379 NETTRAN_DUMMY_12380 NOR2_X1 
XU228 n91 n81 ab_3__11_ NETTRAN_DUMMY_12381 NETTRAN_DUMMY_12382 NOR2_X1 
XU227 n90 n81 ab_3__12_ NETTRAN_DUMMY_12383 NETTRAN_DUMMY_12384 NOR2_X1 
XU226 n89 n81 ab_3__13_ NETTRAN_DUMMY_12385 NETTRAN_DUMMY_12386 NOR2_X1 
XU225 n88 n81 ab_3__14_ NETTRAN_DUMMY_12387 NETTRAN_DUMMY_12388 NOR2_X1 
XU224 n87 n81 ab_3__15_ NETTRAN_DUMMY_12389 NETTRAN_DUMMY_12390 NOR2_X1 
XU223 n86 n81 ab_3__16_ NETTRAN_DUMMY_12391 NETTRAN_DUMMY_12392 NOR2_X1 
XU222 A[3] n85 ab_3__17_ NETTRAN_DUMMY_12393 NETTRAN_DUMMY_12394 NOR2_X1 
XU221 n101 n81 ab_3__1_ NETTRAN_DUMMY_12395 NETTRAN_DUMMY_12396 NOR2_X1 
XU220 n100 n81 ab_3__2_ NETTRAN_DUMMY_12397 NETTRAN_DUMMY_12398 NOR2_X1 
XU219 n99 n81 ab_3__3_ NETTRAN_DUMMY_12399 NETTRAN_DUMMY_12400 NOR2_X1 
XU218 n98 n81 ab_3__4_ NETTRAN_DUMMY_12401 NETTRAN_DUMMY_12402 NOR2_X1 
XU217 n97 n81 ab_3__5_ NETTRAN_DUMMY_12403 NETTRAN_DUMMY_12404 NOR2_X1 
XU216 n96 n81 ab_3__6_ NETTRAN_DUMMY_12405 NETTRAN_DUMMY_12406 NOR2_X1 
XU215 n95 n81 ab_3__7_ NETTRAN_DUMMY_12407 NETTRAN_DUMMY_12408 NOR2_X1 
XU214 n94 n81 ab_3__8_ NETTRAN_DUMMY_12409 NETTRAN_DUMMY_12410 NOR2_X1 
XU213 n93 n81 ab_3__9_ NETTRAN_DUMMY_12411 NETTRAN_DUMMY_12412 NOR2_X1 
XU392 n156 n84 n157 NETTRAN_DUMMY_12413 NETTRAN_DUMMY_12414 NOR2_X1 
XU391 n92 n84 ab_0__10_ NETTRAN_DUMMY_12415 NETTRAN_DUMMY_12416 NOR2_X1 
XU390 n91 n84 ab_0__11_ NETTRAN_DUMMY_12417 NETTRAN_DUMMY_12418 NOR2_X1 
XU389 n90 n84 ab_0__12_ NETTRAN_DUMMY_12419 NETTRAN_DUMMY_12420 NOR2_X1 
XU388 n89 n84 ab_0__13_ NETTRAN_DUMMY_12421 NETTRAN_DUMMY_12422 NOR2_X1 
XU387 n88 n84 ab_0__14_ NETTRAN_DUMMY_12423 NETTRAN_DUMMY_12424 NOR2_X1 
XU386 n87 n84 ab_0__15_ NETTRAN_DUMMY_12425 NETTRAN_DUMMY_12426 NOR2_X1 
XU385 n86 n84 ab_0__16_ NETTRAN_DUMMY_12427 NETTRAN_DUMMY_12428 NOR2_X1 
XU384 A[0] n85 ab_0__17_ NETTRAN_DUMMY_12429 NETTRAN_DUMMY_12430 NOR2_X1 
XU383 n101 n84 ab_0__1_ NETTRAN_DUMMY_12431 NETTRAN_DUMMY_12432 NOR2_X1 
XU382 n100 n84 ab_0__2_ NETTRAN_DUMMY_12433 NETTRAN_DUMMY_12434 NOR2_X1 
XU381 n99 n84 ab_0__3_ NETTRAN_DUMMY_12435 NETTRAN_DUMMY_12436 NOR2_X1 
XU380 n98 n84 ab_0__4_ NETTRAN_DUMMY_12437 NETTRAN_DUMMY_12438 NOR2_X1 
XU379 n97 n84 ab_0__5_ NETTRAN_DUMMY_12439 NETTRAN_DUMMY_12440 NOR2_X1 
XU378 n96 n84 ab_0__6_ NETTRAN_DUMMY_12441 NETTRAN_DUMMY_12442 NOR2_X1 
XU377 n95 n84 ab_0__7_ NETTRAN_DUMMY_12443 NETTRAN_DUMMY_12444 NOR2_X1 
XU376 n94 n84 ab_0__8_ NETTRAN_DUMMY_12445 NETTRAN_DUMMY_12446 NOR2_X1 
XU375 n93 n84 ab_0__9_ NETTRAN_DUMMY_12447 NETTRAN_DUMMY_12448 NOR2_X1 
XU374 n156 n74 ab_10__0_ NETTRAN_DUMMY_12449 NETTRAN_DUMMY_12450 NOR2_X1 
XU373 n92 n74 ab_10__10_ NETTRAN_DUMMY_12451 NETTRAN_DUMMY_12452 NOR2_X1 
XU372 n91 n74 ab_10__11_ NETTRAN_DUMMY_12453 NETTRAN_DUMMY_12454 NOR2_X1 
XU371 n90 n74 ab_10__12_ NETTRAN_DUMMY_12455 NETTRAN_DUMMY_12456 NOR2_X1 
XU370 n89 n74 ab_10__13_ NETTRAN_DUMMY_12457 NETTRAN_DUMMY_12458 NOR2_X1 
XU369 n88 n74 ab_10__14_ NETTRAN_DUMMY_12459 NETTRAN_DUMMY_12460 NOR2_X1 
XU368 n87 n74 ab_10__15_ NETTRAN_DUMMY_12461 NETTRAN_DUMMY_12462 NOR2_X1 
XU367 n86 n74 ab_10__16_ NETTRAN_DUMMY_12463 NETTRAN_DUMMY_12464 NOR2_X1 
XU366 A[10] n85 ab_10__17_ NETTRAN_DUMMY_12465 NETTRAN_DUMMY_12466 NOR2_X1 
XU365 n101 n74 ab_10__1_ NETTRAN_DUMMY_12467 NETTRAN_DUMMY_12468 NOR2_X1 
XU364 n100 n74 ab_10__2_ NETTRAN_DUMMY_12469 NETTRAN_DUMMY_12470 NOR2_X1 
XU363 n99 n74 ab_10__3_ NETTRAN_DUMMY_12471 NETTRAN_DUMMY_12472 NOR2_X1 
XU362 n98 n74 ab_10__4_ NETTRAN_DUMMY_12473 NETTRAN_DUMMY_12474 NOR2_X1 
XU361 n97 n74 ab_10__5_ NETTRAN_DUMMY_12475 NETTRAN_DUMMY_12476 NOR2_X1 
XU360 n96 n74 ab_10__6_ NETTRAN_DUMMY_12477 NETTRAN_DUMMY_12478 NOR2_X1 
XU359 n95 n74 ab_10__7_ NETTRAN_DUMMY_12479 NETTRAN_DUMMY_12480 NOR2_X1 
XU358 n94 n74 ab_10__8_ NETTRAN_DUMMY_12481 NETTRAN_DUMMY_12482 NOR2_X1 
XU357 n93 n74 ab_10__9_ NETTRAN_DUMMY_12483 NETTRAN_DUMMY_12484 NOR2_X1 
XU356 n156 n73 ab_11__0_ NETTRAN_DUMMY_12485 NETTRAN_DUMMY_12486 NOR2_X1 
XU355 n92 n73 ab_11__10_ NETTRAN_DUMMY_12487 NETTRAN_DUMMY_12488 NOR2_X1 
XU354 n91 n73 ab_11__11_ NETTRAN_DUMMY_12489 NETTRAN_DUMMY_12490 NOR2_X1 
XU353 n90 n73 ab_11__12_ NETTRAN_DUMMY_12491 NETTRAN_DUMMY_12492 NOR2_X1 
XU352 n89 n73 ab_11__13_ NETTRAN_DUMMY_12493 NETTRAN_DUMMY_12494 NOR2_X1 
XU351 n88 n73 ab_11__14_ NETTRAN_DUMMY_12495 NETTRAN_DUMMY_12496 NOR2_X1 
XU350 n87 n73 ab_11__15_ NETTRAN_DUMMY_12497 NETTRAN_DUMMY_12498 NOR2_X1 
XU349 n86 n73 ab_11__16_ NETTRAN_DUMMY_12499 NETTRAN_DUMMY_12500 NOR2_X1 
XU348 A[11] n85 ab_11__17_ NETTRAN_DUMMY_12501 NETTRAN_DUMMY_12502 NOR2_X1 
XU347 n101 n73 ab_11__1_ NETTRAN_DUMMY_12503 NETTRAN_DUMMY_12504 NOR2_X1 
XU346 n100 n73 ab_11__2_ NETTRAN_DUMMY_12505 NETTRAN_DUMMY_12506 NOR2_X1 
XU345 n99 n73 ab_11__3_ NETTRAN_DUMMY_12507 NETTRAN_DUMMY_12508 NOR2_X1 
XU344 n98 n73 ab_11__4_ NETTRAN_DUMMY_12509 NETTRAN_DUMMY_12510 NOR2_X1 
XU343 n97 n73 ab_11__5_ NETTRAN_DUMMY_12511 NETTRAN_DUMMY_12512 NOR2_X1 
XU342 n96 n73 ab_11__6_ NETTRAN_DUMMY_12513 NETTRAN_DUMMY_12514 NOR2_X1 
XU341 n95 n73 ab_11__7_ NETTRAN_DUMMY_12515 NETTRAN_DUMMY_12516 NOR2_X1 
XU340 n94 n73 ab_11__8_ NETTRAN_DUMMY_12517 NETTRAN_DUMMY_12518 NOR2_X1 
XU339 n93 n73 ab_11__9_ NETTRAN_DUMMY_12519 NETTRAN_DUMMY_12520 NOR2_X1 
XU338 n156 n72 ab_12__0_ NETTRAN_DUMMY_12521 NETTRAN_DUMMY_12522 NOR2_X1 
XU337 n92 n72 ab_12__10_ NETTRAN_DUMMY_12523 NETTRAN_DUMMY_12524 NOR2_X1 
XU336 n91 n72 ab_12__11_ NETTRAN_DUMMY_12525 NETTRAN_DUMMY_12526 NOR2_X1 
XU335 n90 n72 ab_12__12_ NETTRAN_DUMMY_12527 NETTRAN_DUMMY_12528 NOR2_X1 
XU334 n89 n72 ab_12__13_ NETTRAN_DUMMY_12529 NETTRAN_DUMMY_12530 NOR2_X1 
XU333 n88 n72 ab_12__14_ NETTRAN_DUMMY_12531 NETTRAN_DUMMY_12532 NOR2_X1 
XU332 n87 n72 ab_12__15_ NETTRAN_DUMMY_12533 NETTRAN_DUMMY_12534 NOR2_X1 
XU331 n86 n72 ab_12__16_ NETTRAN_DUMMY_12535 NETTRAN_DUMMY_12536 NOR2_X1 
XU330 A[12] n85 ab_12__17_ NETTRAN_DUMMY_12537 NETTRAN_DUMMY_12538 NOR2_X1 
XU329 n101 n72 ab_12__1_ NETTRAN_DUMMY_12539 NETTRAN_DUMMY_12540 NOR2_X1 
XU328 n100 n72 ab_12__2_ NETTRAN_DUMMY_12541 NETTRAN_DUMMY_12542 NOR2_X1 
XU327 n99 n72 ab_12__3_ NETTRAN_DUMMY_12543 NETTRAN_DUMMY_12544 NOR2_X1 
XU326 n98 n72 ab_12__4_ NETTRAN_DUMMY_12545 NETTRAN_DUMMY_12546 NOR2_X1 
XU325 n97 n72 ab_12__5_ NETTRAN_DUMMY_12547 NETTRAN_DUMMY_12548 NOR2_X1 
XU324 n96 n72 ab_12__6_ NETTRAN_DUMMY_12549 NETTRAN_DUMMY_12550 NOR2_X1 
XU323 n95 n72 ab_12__7_ NETTRAN_DUMMY_12551 NETTRAN_DUMMY_12552 NOR2_X1 
XU322 n94 n72 ab_12__8_ NETTRAN_DUMMY_12553 NETTRAN_DUMMY_12554 NOR2_X1 
XU321 n93 n72 ab_12__9_ NETTRAN_DUMMY_12555 NETTRAN_DUMMY_12556 NOR2_X1 
XU320 n156 n71 ab_13__0_ NETTRAN_DUMMY_12557 NETTRAN_DUMMY_12558 NOR2_X1 
XU319 n92 n71 ab_13__10_ NETTRAN_DUMMY_12559 NETTRAN_DUMMY_12560 NOR2_X1 
XU318 n91 n71 ab_13__11_ NETTRAN_DUMMY_12561 NETTRAN_DUMMY_12562 NOR2_X1 
XU317 n90 n71 ab_13__12_ NETTRAN_DUMMY_12563 NETTRAN_DUMMY_12564 NOR2_X1 
XU316 n89 n71 ab_13__13_ NETTRAN_DUMMY_12565 NETTRAN_DUMMY_12566 NOR2_X1 
XU315 n88 n71 ab_13__14_ NETTRAN_DUMMY_12567 NETTRAN_DUMMY_12568 NOR2_X1 
XU314 n87 n71 ab_13__15_ NETTRAN_DUMMY_12569 NETTRAN_DUMMY_12570 NOR2_X1 
XU313 n86 n71 ab_13__16_ NETTRAN_DUMMY_12571 NETTRAN_DUMMY_12572 NOR2_X1 
XU312 A[13] n85 ab_13__17_ NETTRAN_DUMMY_12573 NETTRAN_DUMMY_12574 NOR2_X1 
XU311 n101 n71 ab_13__1_ NETTRAN_DUMMY_12575 NETTRAN_DUMMY_12576 NOR2_X1 
XU310 n100 n71 ab_13__2_ NETTRAN_DUMMY_12577 NETTRAN_DUMMY_12578 NOR2_X1 
XU309 n99 n71 ab_13__3_ NETTRAN_DUMMY_12579 NETTRAN_DUMMY_12580 NOR2_X1 
XU308 n98 n71 ab_13__4_ NETTRAN_DUMMY_12581 NETTRAN_DUMMY_12582 NOR2_X1 
XU307 n97 n71 ab_13__5_ NETTRAN_DUMMY_12583 NETTRAN_DUMMY_12584 NOR2_X1 
XU306 n96 n71 ab_13__6_ NETTRAN_DUMMY_12585 NETTRAN_DUMMY_12586 NOR2_X1 
XU104 n119 PRODUCT[14] NETTRAN_DUMMY_12587 NETTRAN_DUMMY_12588 BUF_X1 
XU393 n127 PRODUCT[10] NETTRAN_DUMMY_12589 NETTRAN_DUMMY_12590 BUF_X1 
XU394 n129 PRODUCT[9] NETTRAN_DUMMY_12591 NETTRAN_DUMMY_12592 BUF_X1 
XU395 n134 PRODUCT[7] NETTRAN_DUMMY_12593 NETTRAN_DUMMY_12594 BUF_X1 
XU396 n136 PRODUCT[6] NETTRAN_DUMMY_12595 NETTRAN_DUMMY_12596 BUF_X1 
XU397 n138 PRODUCT[5] NETTRAN_DUMMY_12597 NETTRAN_DUMMY_12598 BUF_X1 
XU398 n139 PRODUCT[4] NETTRAN_DUMMY_12599 NETTRAN_DUMMY_12600 BUF_X1 
XU399 n143 PRODUCT[3] NETTRAN_DUMMY_12601 NETTRAN_DUMMY_12602 BUF_X1 
XU400 n144 PRODUCT[2] NETTRAN_DUMMY_12603 NETTRAN_DUMMY_12604 BUF_X1 
XU401 n148 PRODUCT[1] NETTRAN_DUMMY_12605 NETTRAN_DUMMY_12606 BUF_X1 
XU402 n152 PRODUCT[0] NETTRAN_DUMMY_12607 NETTRAN_DUMMY_12608 BUF_X1 
XU403 n102 n155 NETTRAN_DUMMY_12609 NETTRAN_DUMMY_12610 INV_X1 
XU404 n145 n146 NETTRAN_DUMMY_12611 NETTRAN_DUMMY_12612 INV_X1 
XU405 n137 n138 NETTRAN_DUMMY_12613 NETTRAN_DUMMY_12614 INV_X16 
XU406 n140 n141 NETTRAN_DUMMY_12615 NETTRAN_DUMMY_12616 INV_X1 
XU407 n131 n132 NETTRAN_DUMMY_12617 NETTRAN_DUMMY_12618 INV_X1 
XU408 n118 n119 NETTRAN_DUMMY_12619 NETTRAN_DUMMY_12620 INV_X16 
XU409 n117 n114 NETTRAN_DUMMY_12621 NETTRAN_DUMMY_12622 INV_X1 
XU410 n114 PRODUCT[15] NETTRAN_DUMMY_12623 NETTRAN_DUMMY_12624 INV_X32 
XU411 n69 n116 NETTRAN_DUMMY_12625 NETTRAN_DUMMY_12626 INV_X1 
XU412 n116 n117 NETTRAN_DUMMY_12627 NETTRAN_DUMMY_12628 INV_X32 
XU413 A1_12_ n118 NETTRAN_DUMMY_12629 NETTRAN_DUMMY_12630 INV_X32 
XU414 A1_11_ n120 NETTRAN_DUMMY_12631 NETTRAN_DUMMY_12632 INV_X32 
XU415 n120 PRODUCT[13] NETTRAN_DUMMY_12633 NETTRAN_DUMMY_12634 INV_X32 
XU416 A1_10_ n122 NETTRAN_DUMMY_12635 NETTRAN_DUMMY_12636 INV_X32 
XU417 n122 PRODUCT[12] NETTRAN_DUMMY_12637 NETTRAN_DUMMY_12638 INV_X32 
XU418 A1_9_ n124 NETTRAN_DUMMY_12639 NETTRAN_DUMMY_12640 INV_X32 
XU419 n124 n125 NETTRAN_DUMMY_12641 NETTRAN_DUMMY_12642 INV_X32 
XU420 A1_8_ n126 NETTRAN_DUMMY_12643 NETTRAN_DUMMY_12644 INV_X32 
XU421 n126 n127 NETTRAN_DUMMY_12645 NETTRAN_DUMMY_12646 INV_X16 
XU422 A1_7_ n128 NETTRAN_DUMMY_12647 NETTRAN_DUMMY_12648 INV_X32 
XU423 n128 n129 NETTRAN_DUMMY_12649 NETTRAN_DUMMY_12650 INV_X32 
XU424 n132 n130 NETTRAN_DUMMY_12651 NETTRAN_DUMMY_12652 BUF_X1 
XU425 A1_6_ n131 NETTRAN_DUMMY_12653 NETTRAN_DUMMY_12654 INV_X32 
XU426 A1_5_ n133 NETTRAN_DUMMY_12655 NETTRAN_DUMMY_12656 INV_X32 
XU427 n133 n134 NETTRAN_DUMMY_12657 NETTRAN_DUMMY_12658 INV_X32 
XU428 A1_4_ n135 NETTRAN_DUMMY_12659 NETTRAN_DUMMY_12660 INV_X32 
XU429 n135 n136 NETTRAN_DUMMY_12661 NETTRAN_DUMMY_12662 INV_X32 
XU430 A1_3_ n137 NETTRAN_DUMMY_12663 NETTRAN_DUMMY_12664 INV_X32 
XU431 n141 n139 NETTRAN_DUMMY_12665 NETTRAN_DUMMY_12666 BUF_X1 
XU432 A1_2_ n140 NETTRAN_DUMMY_12667 NETTRAN_DUMMY_12668 INV_X32 
XU433 A1_1_ n142 NETTRAN_DUMMY_12669 NETTRAN_DUMMY_12670 INV_X32 
XU434 n142 n143 NETTRAN_DUMMY_12671 NETTRAN_DUMMY_12672 INV_X32 
XU435 n146 n144 NETTRAN_DUMMY_12673 NETTRAN_DUMMY_12674 BUF_X1 
XU436 A1_0_ n145 NETTRAN_DUMMY_12675 NETTRAN_DUMMY_12676 INV_X32 
XU437 n150 n147 NETTRAN_DUMMY_12677 NETTRAN_DUMMY_12678 INV_X1 
XU438 n147 n148 NETTRAN_DUMMY_12679 NETTRAN_DUMMY_12680 INV_X16 
XU439 n158 n149 NETTRAN_DUMMY_12681 NETTRAN_DUMMY_12682 INV_X1 
XU440 n149 n150 NETTRAN_DUMMY_12683 NETTRAN_DUMMY_12684 INV_X32 
XU441 n154 n151 NETTRAN_DUMMY_12685 NETTRAN_DUMMY_12686 INV_X1 
XU442 n151 n152 NETTRAN_DUMMY_12687 NETTRAN_DUMMY_12688 INV_X32 
XU443 n157 n153 NETTRAN_DUMMY_12689 NETTRAN_DUMMY_12690 INV_X1 
XU444 n153 n154 NETTRAN_DUMMY_12691 NETTRAN_DUMMY_12692 INV_X32 
XU445 n155 n156 NETTRAN_DUMMY_12693 NETTRAN_DUMMY_12694 INV_X1 
XU461 n125 PRODUCT[11] NETTRAN_DUMMY_12695 NETTRAN_DUMMY_12696 BUF_X1 
XU462 n130 PRODUCT[8] NETTRAN_DUMMY_12697 NETTRAN_DUMMY_12698 BUF_X1 
XFS_1 VSS NETTRAN_DUMMY_12699 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] PRODUCT[29] 
+ PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] PRODUCT[22] 
+ PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] n49 n61 
+ n60 n59 n58 n57 n56 n55 n54 n53 n52 n51 n50 n41 n40 A2_16_ n39 n68 VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS n70 n48 n67 n47 n66 n46 n65 n45 n64 
+ n44 n63 n43 n62 n37 n42 n36 A1_15_ n38 PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] 
+ PRODUCT[11] PRODUCT[10] PRODUCT[9] PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] 
+ PRODUCT[4] PRODUCT[3] PRODUCT[2] gng_smul_16_18_sadd_37_DW01_add_1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37 p[37] p[36] p[35] p[34] p[33] p[32] p[31] p[30] p[29] 
+ p[28] p[27] p[26] p[25] p[24] p[23] p[22] p[21] p[20] p[19] p[18] p[17] p[16] 
+ p[15] p[14] p[13] p[12] p[11] p[10] p[9] p[8] p[7] p[6] p[5] p[4] p[3] p[2] p[1] 
+ p[0] clk c[36] c[35] c[34] c[33] c[32] c[31] c[30] c[29] c[28] c[27] c[26] c[25] 
+ c[24] c[23] c[22] c[21] c[20] c[19] c[18] c[17] c[16] c[15] c[14] c[13] c[12] 
+ c[11] c[10] c[9] c[8] c[7] c[6] c[5] c[4] c[3] c[2] c[1] c[0] b[17] b[16] b[15] 
+ b[14] b[13] b[12] b[11] b[10] b[9] b[8] b[7] b[6] b[5] b[4] b[3] b[2] b[1] b[0] 
+ a[15] a[14] a[13] a[12] a[11] a[10] a[9] a[8] a[7] a[6] a[5] a[4] a[3] a[2] a[1] 
+ a[0] 
XLOGIC0_X1_U1 LOGIC0_X1_U1_net NETTRAN_DUMMY_12700 NETTRAN_DUMMY_12701 LOGIC0_X1 
XLOGIC0_X1_U2 LOGIC0_X1_U2_net NETTRAN_DUMMY_12702 NETTRAN_DUMMY_12703 LOGIC0_X1 
XLOGIC0_X1_U3 LOGIC0_X1_U3_net NETTRAN_DUMMY_12704 NETTRAN_DUMMY_12705 LOGIC0_X1 
XLOGIC0_X1_U4 LOGIC0_X1_U4_net NETTRAN_DUMMY_12706 NETTRAN_DUMMY_12707 LOGIC0_X1 
Xprod_reg_30_ N301 n2_G3B1I6 prod[30] NETTRAN_DUMMY_12708 NETTRAN_DUMMY_12709 NETTRAN_DUMMY_12710 DFF_X1 
Xprod_reg_31_ N310 n2_G3B1I6 prod[31] NETTRAN_DUMMY_12711 NETTRAN_DUMMY_12712 NETTRAN_DUMMY_12713 DFF_X1 
Xprod_reg_32_ N320 n2_G3B1I2 prod[32] NETTRAN_DUMMY_12714 NETTRAN_DUMMY_12715 NETTRAN_DUMMY_12716 DFF_X1 
Xprod_reg_33_ N33 n2_G3B1I2 prod[33] NETTRAN_DUMMY_12717 NETTRAN_DUMMY_12718 NETTRAN_DUMMY_12719 DFF_X1 
Xc_reg_reg_0_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[0] NETTRAN_DUMMY_12720 NETTRAN_DUMMY_12721 
+ NETTRAN_DUMMY_12722 DFF_X1 
Xc_reg_reg_1_ LOGIC0_X1_U4_net n3 c_reg[1] NETTRAN_DUMMY_12723 NETTRAN_DUMMY_12724 
+ NETTRAN_DUMMY_12725 DFF_X1 
Xc_reg_reg_2_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[2] NETTRAN_DUMMY_12726 NETTRAN_DUMMY_12727 
+ NETTRAN_DUMMY_12728 DFF_X1 
Xc_reg_reg_3_ LOGIC0_X1_U4_net n3 c_reg[3] NETTRAN_DUMMY_12729 NETTRAN_DUMMY_12730 
+ NETTRAN_DUMMY_12731 DFF_X1 
Xc_reg_reg_4_ LOGIC0_X1_U4_net n3 c_reg[4] NETTRAN_DUMMY_12732 NETTRAN_DUMMY_12733 
+ NETTRAN_DUMMY_12734 DFF_X1 
Xc_reg_reg_5_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[5] NETTRAN_DUMMY_12735 NETTRAN_DUMMY_12736 
+ NETTRAN_DUMMY_12737 DFF_X1 
Xc_reg_reg_6_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[6] NETTRAN_DUMMY_12738 NETTRAN_DUMMY_12739 
+ NETTRAN_DUMMY_12740 DFF_X1 
Xc_reg_reg_7_ LOGIC0_X1_U4_net n3_G3B1I4 c_reg[7] NETTRAN_DUMMY_12741 NETTRAN_DUMMY_12742 
+ NETTRAN_DUMMY_12743 DFF_X1 
Xc_reg_reg_8_ LOGIC0_X1_U3_net n3_G3B1I4 c_reg[8] NETTRAN_DUMMY_12744 NETTRAN_DUMMY_12745 
+ NETTRAN_DUMMY_12746 DFF_X1 
Xc_reg_reg_9_ LOGIC0_X1_U4_net n3_G3B1I4 c_reg[9] NETTRAN_DUMMY_12747 NETTRAN_DUMMY_12748 
+ NETTRAN_DUMMY_12749 DFF_X1 
Xc_reg_reg_10_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[10] NETTRAN_DUMMY_12750 NETTRAN_DUMMY_12751 
+ NETTRAN_DUMMY_12752 DFF_X1 
Xc_reg_reg_11_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[11] NETTRAN_DUMMY_12753 NETTRAN_DUMMY_12754 
+ NETTRAN_DUMMY_12755 DFF_X1 
Xc_reg_reg_12_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[12] NETTRAN_DUMMY_12756 NETTRAN_DUMMY_12757 
+ NETTRAN_DUMMY_12758 DFF_X1 
Xc_reg_reg_13_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[13] NETTRAN_DUMMY_12759 NETTRAN_DUMMY_12760 
+ NETTRAN_DUMMY_12761 DFF_X1 
Xc_reg_reg_14_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[14] NETTRAN_DUMMY_12762 NETTRAN_DUMMY_12763 
+ NETTRAN_DUMMY_12764 DFF_X1 
Xc_reg_reg_15_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[15] NETTRAN_DUMMY_12765 NETTRAN_DUMMY_12766 
+ NETTRAN_DUMMY_12767 DFF_X1 
Xc_reg_reg_16_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[16] NETTRAN_DUMMY_12768 NETTRAN_DUMMY_12769 
+ NETTRAN_DUMMY_12770 DFF_X1 
Xc_reg_reg_17_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[17] NETTRAN_DUMMY_12771 NETTRAN_DUMMY_12772 
+ NETTRAN_DUMMY_12773 DFF_X1 
Xc_reg_reg_18_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[18] NETTRAN_DUMMY_12774 NETTRAN_DUMMY_12775 
+ NETTRAN_DUMMY_12776 DFF_X1 
Xc_reg_reg_19_ c[19] n1_G3B1I6 c_reg[19] NETTRAN_DUMMY_12777 NETTRAN_DUMMY_12778 
+ NETTRAN_DUMMY_12779 DFF_X1 
Xc_reg_reg_20_ c[20] n1_G3B1I3 c_reg[20] NETTRAN_DUMMY_12780 NETTRAN_DUMMY_12781 
+ NETTRAN_DUMMY_12782 DFF_X1 
Xc_reg_reg_21_ c[21] n1_G3B1I3 c_reg[21] NETTRAN_DUMMY_12783 NETTRAN_DUMMY_12784 
+ NETTRAN_DUMMY_12785 DFF_X1 
Xc_reg_reg_22_ c[22] n1_G3B1I3 c_reg[22] NETTRAN_DUMMY_12786 NETTRAN_DUMMY_12787 
+ NETTRAN_DUMMY_12788 DFF_X1 
Xc_reg_reg_23_ c[23] n1_G3B1I3 c_reg[23] NETTRAN_DUMMY_12789 NETTRAN_DUMMY_12790 
+ NETTRAN_DUMMY_12791 DFF_X1 
Xc_reg_reg_24_ c[24] n2_G3B1I3 c_reg[24] NETTRAN_DUMMY_12792 NETTRAN_DUMMY_12793 
+ NETTRAN_DUMMY_12794 DFF_X1 
Xc_reg_reg_25_ c[25] n2_G3B1I3 c_reg[25] NETTRAN_DUMMY_12795 NETTRAN_DUMMY_12796 
+ NETTRAN_DUMMY_12797 DFF_X1 
Xc_reg_reg_26_ c[26] n2_G3B1I3 c_reg[26] NETTRAN_DUMMY_12798 NETTRAN_DUMMY_12799 
+ NETTRAN_DUMMY_12800 DFF_X1 
Xc_reg_reg_27_ c[27] n2_G3B1I3 c_reg[27] NETTRAN_DUMMY_12801 NETTRAN_DUMMY_12802 
+ NETTRAN_DUMMY_12803 DFF_X1 
Xc_reg_reg_28_ c[28] n2_G3B1I3 c_reg[28] NETTRAN_DUMMY_12804 NETTRAN_DUMMY_12805 
+ NETTRAN_DUMMY_12806 DFF_X1 
Xc_reg_reg_29_ c[29] n2_G3B1I3 c_reg[29] NETTRAN_DUMMY_12807 NETTRAN_DUMMY_12808 
+ NETTRAN_DUMMY_12809 DFF_X1 
Xc_reg_reg_30_ c[30] n2_G3B1I3 c_reg[30] NETTRAN_DUMMY_12810 NETTRAN_DUMMY_12811 
+ NETTRAN_DUMMY_12812 DFF_X1 
Xc_reg_reg_31_ c[31] n2_G3B1I4 c_reg[31] NETTRAN_DUMMY_12813 NETTRAN_DUMMY_12814 
+ NETTRAN_DUMMY_12815 DFF_X1 
Xc_reg_reg_32_ c[32] n2_G3B1I4 c_reg[32] NETTRAN_DUMMY_12816 NETTRAN_DUMMY_12817 
+ NETTRAN_DUMMY_12818 DFF_X1 
Xc_reg_reg_33_ c[33] n2_G3B1I4 c_reg[33] NETTRAN_DUMMY_12819 NETTRAN_DUMMY_12820 
+ NETTRAN_DUMMY_12821 DFF_X1 
Xc_reg_reg_34_ c[34] n2_G3B1I2 c_reg[34] NETTRAN_DUMMY_12822 NETTRAN_DUMMY_12823 
+ NETTRAN_DUMMY_12824 DFF_X1 
Xc_reg_reg_35_ c[35] n2_G3B1I2 c_reg[35] NETTRAN_DUMMY_12825 NETTRAN_DUMMY_12826 
+ NETTRAN_DUMMY_12827 DFF_X1 
Xc_reg_reg_36_ c[36] n2_G3B1I2 c_reg[36] NETTRAN_DUMMY_12828 NETTRAN_DUMMY_12829 
+ NETTRAN_DUMMY_12830 DFF_X1 
Xb_reg_reg_0_ b[0] n2_G3B1I1 b_reg[0] NETTRAN_DUMMY_12831 NETTRAN_DUMMY_12832 NETTRAN_DUMMY_12833 DFF_X1 
Xb_reg_reg_1_ b[1] n2_G3B1I1 b_reg[1] NETTRAN_DUMMY_12834 NETTRAN_DUMMY_12835 NETTRAN_DUMMY_12836 DFF_X1 
Xb_reg_reg_2_ b[2] n1_G3B1I6 b_reg[2] NETTRAN_DUMMY_12837 NETTRAN_DUMMY_12838 NETTRAN_DUMMY_12839 DFF_X1 
Xb_reg_reg_3_ b[3] n1_G3B1I6 b_reg[3] NETTRAN_DUMMY_12840 NETTRAN_DUMMY_12841 NETTRAN_DUMMY_12842 DFF_X1 
Xb_reg_reg_4_ b[4] n1_G3B1I2 b_reg[4] NETTRAN_DUMMY_12843 NETTRAN_DUMMY_12844 NETTRAN_DUMMY_12845 DFF_X1 
Xb_reg_reg_5_ b[5] n1_G3B1I2 b_reg[5] NETTRAN_DUMMY_12846 NETTRAN_DUMMY_12847 NETTRAN_DUMMY_12848 DFF_X1 
Xb_reg_reg_6_ b[6] n1_G3B1I2 b_reg[6] NETTRAN_DUMMY_12849 NETTRAN_DUMMY_12850 NETTRAN_DUMMY_12851 DFF_X1 
Xb_reg_reg_7_ b[7] n1_G3B1I3 b_reg[7] NETTRAN_DUMMY_12852 NETTRAN_DUMMY_12853 NETTRAN_DUMMY_12854 DFF_X1 
Xb_reg_reg_8_ b[8] n1_G3B1I4 b_reg[8] NETTRAN_DUMMY_12855 NETTRAN_DUMMY_12856 NETTRAN_DUMMY_12857 DFF_X1 
Xb_reg_reg_9_ b[9] n1_G3B1I4 b_reg[9] NETTRAN_DUMMY_12858 NETTRAN_DUMMY_12859 NETTRAN_DUMMY_12860 DFF_X1 
Xb_reg_reg_10_ b[10] n2_G3B1I1 b_reg[10] NETTRAN_DUMMY_12861 NETTRAN_DUMMY_12862 
+ NETTRAN_DUMMY_12863 DFF_X1 
Xb_reg_reg_11_ b[11] n2_G3B1I6 b_reg[11] NETTRAN_DUMMY_12864 NETTRAN_DUMMY_12865 
+ NETTRAN_DUMMY_12866 DFF_X1 
Xb_reg_reg_12_ b[12] n2_G3B1I1 b_reg[12] NETTRAN_DUMMY_12867 NETTRAN_DUMMY_12868 
+ NETTRAN_DUMMY_12869 DFF_X1 
Xb_reg_reg_13_ b[13] n2_G3B1I6 b_reg[13] NETTRAN_DUMMY_12870 NETTRAN_DUMMY_12871 
+ NETTRAN_DUMMY_12872 DFF_X1 
Xb_reg_reg_14_ b[14] n2_G3B1I1 b_reg[14] NETTRAN_DUMMY_12873 NETTRAN_DUMMY_12874 
+ NETTRAN_DUMMY_12875 DFF_X1 
Xb_reg_reg_15_ b[15] n2_G3B1I1 b_reg[15] NETTRAN_DUMMY_12876 NETTRAN_DUMMY_12877 
+ NETTRAN_DUMMY_12878 DFF_X1 
Xb_reg_reg_16_ b[16] n2_G3B1I1 b_reg[16] NETTRAN_DUMMY_12879 NETTRAN_DUMMY_12880 
+ NETTRAN_DUMMY_12881 DFF_X1 
Xb_reg_reg_17_ LOGIC0_X1_U2_net n1_G3B1I2 b_reg[17] NETTRAN_DUMMY_12882 NETTRAN_DUMMY_12883 
+ NETTRAN_DUMMY_12884 DFF_X1 
Xa_reg_reg_0_ a[0] n1_G3B1I6 a_reg[0] NETTRAN_DUMMY_12885 NETTRAN_DUMMY_12886 NETTRAN_DUMMY_12887 DFF_X1 
Xa_reg_reg_1_ a[1] n1_G3B1I6 a_reg[1] NETTRAN_DUMMY_12888 NETTRAN_DUMMY_12889 NETTRAN_DUMMY_12890 DFF_X1 
Xa_reg_reg_2_ a[2] n1_G3B1I2 a_reg[2] NETTRAN_DUMMY_12891 NETTRAN_DUMMY_12892 NETTRAN_DUMMY_12893 DFF_X1 
Xa_reg_reg_3_ a[3] n1_G3B1I6 a_reg[3] NETTRAN_DUMMY_12894 NETTRAN_DUMMY_12895 NETTRAN_DUMMY_12896 DFF_X1 
Xa_reg_reg_4_ a[4] n1_G3B1I1 a_reg[4] NETTRAN_DUMMY_12897 NETTRAN_DUMMY_12898 NETTRAN_DUMMY_12899 DFF_X1 
Xa_reg_reg_5_ a[5] n1_G3B1I2 a_reg[5] NETTRAN_DUMMY_12900 NETTRAN_DUMMY_12901 NETTRAN_DUMMY_12902 DFF_X1 
Xa_reg_reg_6_ a[6] n1_G3B1I1 a_reg[6] NETTRAN_DUMMY_12903 NETTRAN_DUMMY_12904 NETTRAN_DUMMY_12905 DFF_X1 
Xa_reg_reg_7_ a[7] n1_G3B1I1 a_reg[7] NETTRAN_DUMMY_12906 NETTRAN_DUMMY_12907 NETTRAN_DUMMY_12908 DFF_X1 
Xa_reg_reg_8_ a[8] n1_G3B1I1 a_reg[8] NETTRAN_DUMMY_12909 NETTRAN_DUMMY_12910 NETTRAN_DUMMY_12911 DFF_X1 
Xa_reg_reg_9_ a[9] n2 a_reg[9] NETTRAN_DUMMY_12912 NETTRAN_DUMMY_12913 NETTRAN_DUMMY_12914 DFF_X1 
Xa_reg_reg_10_ a[10] n1_G3B1I4 a_reg[10] NETTRAN_DUMMY_12915 NETTRAN_DUMMY_12916 
+ NETTRAN_DUMMY_12917 DFF_X1 
Xa_reg_reg_11_ a[11] n1_G3B1I4 a_reg[11] NETTRAN_DUMMY_12918 NETTRAN_DUMMY_12919 
+ NETTRAN_DUMMY_12920 DFF_X1 
Xa_reg_reg_12_ a[12] n1_G3B1I4 a_reg[12] NETTRAN_DUMMY_12921 NETTRAN_DUMMY_12922 
+ NETTRAN_DUMMY_12923 DFF_X1 
Xa_reg_reg_13_ a[13] n1_G3B1I4 a_reg[13] NETTRAN_DUMMY_12924 NETTRAN_DUMMY_12925 
+ NETTRAN_DUMMY_12926 DFF_X1 
Xa_reg_reg_14_ a[14] n1_G3B1I4 a_reg[14] NETTRAN_DUMMY_12927 NETTRAN_DUMMY_12928 
+ NETTRAN_DUMMY_12929 DFF_X1 
Xa_reg_reg_15_ LOGIC0_X1_U2_net n1_G3B1I1 a_reg[15] NETTRAN_DUMMY_12930 NETTRAN_DUMMY_12931 
+ NETTRAN_DUMMY_12932 DFF_X1 
Xresult_reg_20_ sum[20] n1_G3B1I3 n119 NETTRAN_DUMMY_12933 NETTRAN_DUMMY_12934 NETTRAN_DUMMY_12935 DFF_X1 
Xresult_reg_21_ sum[21] n1_G3B1I3 n120 NETTRAN_DUMMY_12936 NETTRAN_DUMMY_12937 NETTRAN_DUMMY_12938 DFF_X1 
Xresult_reg_22_ sum[22] n1_G3B1I4 n121 NETTRAN_DUMMY_12939 NETTRAN_DUMMY_12940 NETTRAN_DUMMY_12941 DFF_X1 
Xresult_reg_23_ sum[23] n1_G3B1I4 n122 NETTRAN_DUMMY_12942 NETTRAN_DUMMY_12943 NETTRAN_DUMMY_12944 DFF_X1 
Xresult_reg_24_ sum[24] n2_G3B1I2 n123 NETTRAN_DUMMY_12945 NETTRAN_DUMMY_12946 NETTRAN_DUMMY_12947 DFF_X1 
Xresult_reg_25_ n124 n2_G3B1I3 n111 NETTRAN_DUMMY_12948 NETTRAN_DUMMY_12949 NETTRAN_DUMMY_12950 DFF_X1 
Xresult_reg_26_ sum[26] n2_G3B1I5 n112 NETTRAN_DUMMY_12951 NETTRAN_DUMMY_12952 NETTRAN_DUMMY_12953 DFF_X1 
Xresult_reg_27_ sum[27] n2_G3B1I5 n113 NETTRAN_DUMMY_12954 NETTRAN_DUMMY_12955 NETTRAN_DUMMY_12956 DFF_X1 
Xresult_reg_28_ sum[28] n2_G3B1I5 n114 NETTRAN_DUMMY_12957 NETTRAN_DUMMY_12958 NETTRAN_DUMMY_12959 DFF_X1 
Xresult_reg_29_ sum[29] n2_G3B1I5 n115 NETTRAN_DUMMY_12960 NETTRAN_DUMMY_12961 NETTRAN_DUMMY_12962 DFF_X1 
Xresult_reg_30_ sum[30] n2_G3B1I5 n116 NETTRAN_DUMMY_12963 NETTRAN_DUMMY_12964 NETTRAN_DUMMY_12965 DFF_X1 
Xresult_reg_31_ sum[31] n2_G3B1I4 n117 NETTRAN_DUMMY_12966 NETTRAN_DUMMY_12967 NETTRAN_DUMMY_12968 DFF_X1 
Xresult_reg_32_ sum[32] n2_G3B1I4 n118 NETTRAN_DUMMY_12969 NETTRAN_DUMMY_12970 NETTRAN_DUMMY_12971 DFF_X1 
Xresult_reg_33_ sum[33] n2_G3B1I4 n106 NETTRAN_DUMMY_12972 NETTRAN_DUMMY_12973 NETTRAN_DUMMY_12974 DFF_X1 
Xresult_reg_34_ sum[34] n2_G3B1I4 n107 NETTRAN_DUMMY_12975 NETTRAN_DUMMY_12976 NETTRAN_DUMMY_12977 DFF_X1 
Xresult_reg_35_ sum[35] n2_G3B1I2 n108 NETTRAN_DUMMY_12978 NETTRAN_DUMMY_12979 NETTRAN_DUMMY_12980 DFF_X1 
Xresult_reg_36_ sum[36] n2_G3B1I2 n109 NETTRAN_DUMMY_12981 NETTRAN_DUMMY_12982 NETTRAN_DUMMY_12983 DFF_X1 
Xresult_reg_37_ sum[37] n2_G3B1I6 n110 NETTRAN_DUMMY_12984 NETTRAN_DUMMY_12985 NETTRAN_DUMMY_12986 DFF_X1 
Xprod_reg_0_ N0 n3_G3B1I5 prod[0] NETTRAN_DUMMY_12987 NETTRAN_DUMMY_12988 NETTRAN_DUMMY_12989 DFF_X1 
Xprod_reg_1_ N1000 n3_G3B1I5 prod[1] NETTRAN_DUMMY_12990 NETTRAN_DUMMY_12991 NETTRAN_DUMMY_12992 DFF_X1 
Xprod_reg_2_ N200 n3_G3B1I5 prod[2] NETTRAN_DUMMY_12993 NETTRAN_DUMMY_12994 NETTRAN_DUMMY_12995 DFF_X1 
Xprod_reg_3_ N300 n3_G3B1I5 prod[3] NETTRAN_DUMMY_12996 NETTRAN_DUMMY_12997 NETTRAN_DUMMY_12998 DFF_X1 
Xprod_reg_4_ N4 n3_G3B1I5 prod[4] NETTRAN_DUMMY_12999 NETTRAN_DUMMY_13000 NETTRAN_DUMMY_13001 DFF_X1 
Xprod_reg_5_ N5 n3_G3B1I3 prod[5] NETTRAN_DUMMY_13002 NETTRAN_DUMMY_13003 NETTRAN_DUMMY_13004 DFF_X1 
Xprod_reg_6_ N6 n3_G3B1I3 prod[6] NETTRAN_DUMMY_13005 NETTRAN_DUMMY_13006 NETTRAN_DUMMY_13007 DFF_X1 
Xprod_reg_7_ N7 n3_G3B1I4 prod[7] NETTRAN_DUMMY_13008 NETTRAN_DUMMY_13009 NETTRAN_DUMMY_13010 DFF_X1 
Xprod_reg_8_ N8 n3_G3B1I4 prod[8] NETTRAN_DUMMY_13011 NETTRAN_DUMMY_13012 NETTRAN_DUMMY_13013 DFF_X1 
Xprod_reg_9_ N9 n3_G3B1I4 prod[9] NETTRAN_DUMMY_13014 NETTRAN_DUMMY_13015 NETTRAN_DUMMY_13016 DFF_X1 
Xprod_reg_10_ N102 n3_G3B1I3 prod[10] NETTRAN_DUMMY_13017 NETTRAN_DUMMY_13018 NETTRAN_DUMMY_13019 DFF_X1 
Xprod_reg_11_ N11 n3_G3B1I2 prod[11] NETTRAN_DUMMY_13020 NETTRAN_DUMMY_13021 NETTRAN_DUMMY_13022 DFF_X1 
Xprod_reg_12_ N12 n3_G3B1I2 prod[12] NETTRAN_DUMMY_13023 NETTRAN_DUMMY_13024 NETTRAN_DUMMY_13025 DFF_X1 
Xprod_reg_13_ N13 n3_G3B1I2 prod[13] NETTRAN_DUMMY_13026 NETTRAN_DUMMY_13027 NETTRAN_DUMMY_13028 DFF_X1 
Xprod_reg_14_ N14 n3_G3B1I2 prod[14] NETTRAN_DUMMY_13029 NETTRAN_DUMMY_13030 NETTRAN_DUMMY_13031 DFF_X1 
Xprod_reg_15_ N15 n3_G3B1I2 prod[15] NETTRAN_DUMMY_13032 NETTRAN_DUMMY_13033 NETTRAN_DUMMY_13034 DFF_X1 
Xprod_reg_16_ N16 n1_G3B1I5 prod[16] NETTRAN_DUMMY_13035 NETTRAN_DUMMY_13036 NETTRAN_DUMMY_13037 DFF_X1 
Xprod_reg_17_ N17 n1_G3B1I5 prod[17] NETTRAN_DUMMY_13038 NETTRAN_DUMMY_13039 NETTRAN_DUMMY_13040 DFF_X1 
Xprod_reg_18_ N18 n1_G3B1I5 prod[18] NETTRAN_DUMMY_13041 NETTRAN_DUMMY_13042 NETTRAN_DUMMY_13043 DFF_X1 
Xprod_reg_19_ N19 n1_G3B1I6 prod[19] NETTRAN_DUMMY_13044 NETTRAN_DUMMY_13045 NETTRAN_DUMMY_13046 DFF_X1 
Xprod_reg_20_ N201 n1_G3B1I6 prod[20] NETTRAN_DUMMY_13047 NETTRAN_DUMMY_13048 NETTRAN_DUMMY_13049 DFF_X1 
Xprod_reg_21_ N21 n1_G3B1I3 prod[21] NETTRAN_DUMMY_13050 NETTRAN_DUMMY_13051 NETTRAN_DUMMY_13052 DFF_X1 
Xprod_reg_22_ N22 n1_G3B1I3 prod[22] NETTRAN_DUMMY_13053 NETTRAN_DUMMY_13054 NETTRAN_DUMMY_13055 DFF_X1 
Xprod_reg_23_ N23 n1_G3B1I4 prod[23] NETTRAN_DUMMY_13056 NETTRAN_DUMMY_13057 NETTRAN_DUMMY_13058 DFF_X1 
Xprod_reg_24_ N24 n2_G3B1I1 prod[24] NETTRAN_DUMMY_13059 NETTRAN_DUMMY_13060 NETTRAN_DUMMY_13061 DFF_X1 
Xprod_reg_25_ N25 n2_G3B1I6 prod[25] NETTRAN_DUMMY_13062 NETTRAN_DUMMY_13063 NETTRAN_DUMMY_13064 DFF_X1 
Xprod_reg_26_ N26 n2_G3B1I6 prod[26] NETTRAN_DUMMY_13065 NETTRAN_DUMMY_13066 NETTRAN_DUMMY_13067 DFF_X1 
Xprod_reg_27_ N27 n2_G3B1I6 prod[27] NETTRAN_DUMMY_13068 NETTRAN_DUMMY_13069 NETTRAN_DUMMY_13070 DFF_X1 
Xprod_reg_28_ N28 n2_G3B1I6 prod[28] NETTRAN_DUMMY_13071 NETTRAN_DUMMY_13072 NETTRAN_DUMMY_13073 DFF_X1 
Xprod_reg_29_ N290 n2_G3B1I6 prod[29] NETTRAN_DUMMY_13074 NETTRAN_DUMMY_13075 NETTRAN_DUMMY_13076 DFF_X1 
XU1 clk n1 NETTRAN_DUMMY_13077 NETTRAN_DUMMY_13078 BUF_X32 
XU2 clk n2 NETTRAN_DUMMY_13079 NETTRAN_DUMMY_13080 BUF_X32 
XU3 clk n3 NETTRAN_DUMMY_13081 NETTRAN_DUMMY_13082 BUF_X32 
XCLKBUF_X1_G3B1I61 n1 n1_G3B1I6 NETTRAN_DUMMY_13083 NETTRAN_DUMMY_13084 CLKBUF_X2 
XCLKBUF_X1_G3B1I52 n1 n1_G3B1I5 NETTRAN_DUMMY_13085 NETTRAN_DUMMY_13086 CLKBUF_X2 
XCLKBUF_X1_G3B1I32 n1 n1_G3B1I3 NETTRAN_DUMMY_13087 NETTRAN_DUMMY_13088 CLKBUF_X2 
XCLKBUF_X1_G3B1I22 n1 n1_G3B1I2 NETTRAN_DUMMY_13089 NETTRAN_DUMMY_13090 CLKBUF_X2 
XCLKBUF_X1_G3B1I12 n1 n1_G3B1I1 NETTRAN_DUMMY_13091 NETTRAN_DUMMY_13092 CLKBUF_X2 
XCLKBUF_X1_G3B1I5 n3 n3_G3B1I5 NETTRAN_DUMMY_13093 NETTRAN_DUMMY_13094 CLKBUF_X2 
XCLKBUF_X1_G3B1I4 n3 n3_G3B1I4 NETTRAN_DUMMY_13095 NETTRAN_DUMMY_13096 CLKBUF_X2 
XCLKBUF_X1_G3B1I3 n3 n3_G3B1I3 NETTRAN_DUMMY_13097 NETTRAN_DUMMY_13098 CLKBUF_X2 
XCLKBUF_X1_G3B1I2 n3 n3_G3B1I2 NETTRAN_DUMMY_13099 NETTRAN_DUMMY_13100 CLKBUF_X2 
XCLKBUF_X1_G3B1I6 n2 n2_G3B1I6 NETTRAN_DUMMY_13101 NETTRAN_DUMMY_13102 CLKBUF_X2 
XCLKBUF_X1_G3B1I51 n2 n2_G3B1I5 NETTRAN_DUMMY_13103 NETTRAN_DUMMY_13104 CLKBUF_X2 
XCLKBUF_X1_G3B1I41 n2 n2_G3B1I4 NETTRAN_DUMMY_13105 NETTRAN_DUMMY_13106 CLKBUF_X2 
XCLKBUF_X1_G3B1I31 n2 n2_G3B1I3 NETTRAN_DUMMY_13107 NETTRAN_DUMMY_13108 CLKBUF_X2 
XCLKBUF_X1_G3B1I21 n2 n2_G3B1I2 NETTRAN_DUMMY_13109 NETTRAN_DUMMY_13110 CLKBUF_X2 
XCLKBUF_X1_G3B1I11 n2 n2_G3B1I1 NETTRAN_DUMMY_13111 NETTRAN_DUMMY_13112 CLKBUF_X2 
XCLKBUF_X1_G3B1I42 n1 n1_G3B1I4 NETTRAN_DUMMY_13113 NETTRAN_DUMMY_13114 CLKBUF_X2 
XU4 n31 n330 NETTRAN_DUMMY_13115 NETTRAN_DUMMY_13116 INV_X16 
XU5 b_reg[17] n29 NETTRAN_DUMMY_13117 NETTRAN_DUMMY_13118 INV_X16 
XU6 a_reg[15] n32 NETTRAN_DUMMY_13119 NETTRAN_DUMMY_13120 INV_X1 
XU7 n29 n302 NETTRAN_DUMMY_13121 NETTRAN_DUMMY_13122 INV_X1 
XU8 n32 n31 NETTRAN_DUMMY_13123 NETTRAN_DUMMY_13124 CLKBUF_X1 
XU9 n110 n34 NETTRAN_DUMMY_13125 NETTRAN_DUMMY_13126 CLKBUF_X1 
XU10 n36 n35 NETTRAN_DUMMY_13127 NETTRAN_DUMMY_13128 CLKBUF_X1 
XU11 n34 n36 NETTRAN_DUMMY_13129 NETTRAN_DUMMY_13130 INV_X32 
XU12 n35 p[37] NETTRAN_DUMMY_13131 NETTRAN_DUMMY_13132 INV_X32 
XU13 n109 n38 NETTRAN_DUMMY_13133 NETTRAN_DUMMY_13134 CLKBUF_X1 
XU14 n40 n39 NETTRAN_DUMMY_13135 NETTRAN_DUMMY_13136 CLKBUF_X1 
XU15 n38 n40 NETTRAN_DUMMY_13137 NETTRAN_DUMMY_13138 INV_X32 
XU16 n39 p[36] NETTRAN_DUMMY_13139 NETTRAN_DUMMY_13140 INV_X32 
XU17 n108 n42 NETTRAN_DUMMY_13141 NETTRAN_DUMMY_13142 CLKBUF_X1 
XU18 n44 n43 NETTRAN_DUMMY_13143 NETTRAN_DUMMY_13144 CLKBUF_X1 
XU19 n42 n44 NETTRAN_DUMMY_13145 NETTRAN_DUMMY_13146 INV_X32 
XU20 n43 p[35] NETTRAN_DUMMY_13147 NETTRAN_DUMMY_13148 INV_X32 
XU21 n107 n46 NETTRAN_DUMMY_13149 NETTRAN_DUMMY_13150 CLKBUF_X1 
XU22 n48 n47 NETTRAN_DUMMY_13151 NETTRAN_DUMMY_13152 CLKBUF_X1 
XU23 n46 n48 NETTRAN_DUMMY_13153 NETTRAN_DUMMY_13154 INV_X32 
XU24 n47 p[34] NETTRAN_DUMMY_13155 NETTRAN_DUMMY_13156 INV_X32 
XU25 n106 n50 NETTRAN_DUMMY_13157 NETTRAN_DUMMY_13158 CLKBUF_X1 
XU26 n52 n51 NETTRAN_DUMMY_13159 NETTRAN_DUMMY_13160 CLKBUF_X1 
XU27 n50 n52 NETTRAN_DUMMY_13161 NETTRAN_DUMMY_13162 INV_X32 
XU28 n51 p[33] NETTRAN_DUMMY_13163 NETTRAN_DUMMY_13164 INV_X32 
XU29 n118 n54 NETTRAN_DUMMY_13165 NETTRAN_DUMMY_13166 CLKBUF_X1 
XU30 n56 n55 NETTRAN_DUMMY_13167 NETTRAN_DUMMY_13168 CLKBUF_X1 
XU31 n54 n56 NETTRAN_DUMMY_13169 NETTRAN_DUMMY_13170 INV_X32 
XU32 n55 p[32] NETTRAN_DUMMY_13171 NETTRAN_DUMMY_13172 INV_X32 
XU33 n117 n58 NETTRAN_DUMMY_13173 NETTRAN_DUMMY_13174 CLKBUF_X1 
XU34 n60 n59 NETTRAN_DUMMY_13175 NETTRAN_DUMMY_13176 CLKBUF_X1 
XU35 n58 n60 NETTRAN_DUMMY_13177 NETTRAN_DUMMY_13178 INV_X32 
XU36 n59 p[31] NETTRAN_DUMMY_13179 NETTRAN_DUMMY_13180 INV_X32 
XU37 n116 n62 NETTRAN_DUMMY_13181 NETTRAN_DUMMY_13182 CLKBUF_X1 
XU38 n64 n63 NETTRAN_DUMMY_13183 NETTRAN_DUMMY_13184 CLKBUF_X1 
XU39 n62 n64 NETTRAN_DUMMY_13185 NETTRAN_DUMMY_13186 INV_X32 
XU40 n63 p[30] NETTRAN_DUMMY_13187 NETTRAN_DUMMY_13188 INV_X32 
XU41 n115 n66 NETTRAN_DUMMY_13189 NETTRAN_DUMMY_13190 CLKBUF_X1 
XU42 n68 n67 NETTRAN_DUMMY_13191 NETTRAN_DUMMY_13192 CLKBUF_X1 
XU43 n66 n68 NETTRAN_DUMMY_13193 NETTRAN_DUMMY_13194 INV_X32 
XU44 n67 p[29] NETTRAN_DUMMY_13195 NETTRAN_DUMMY_13196 INV_X32 
XU45 n114 n70 NETTRAN_DUMMY_13197 NETTRAN_DUMMY_13198 CLKBUF_X1 
XU46 n72 n71 NETTRAN_DUMMY_13199 NETTRAN_DUMMY_13200 CLKBUF_X1 
XU47 n70 n72 NETTRAN_DUMMY_13201 NETTRAN_DUMMY_13202 INV_X32 
XU48 n71 p[28] NETTRAN_DUMMY_13203 NETTRAN_DUMMY_13204 INV_X32 
XU49 n113 n74 NETTRAN_DUMMY_13205 NETTRAN_DUMMY_13206 CLKBUF_X1 
XU50 n76 n75 NETTRAN_DUMMY_13207 NETTRAN_DUMMY_13208 CLKBUF_X1 
XU51 n74 n76 NETTRAN_DUMMY_13209 NETTRAN_DUMMY_13210 INV_X32 
XU52 n75 p[27] NETTRAN_DUMMY_13211 NETTRAN_DUMMY_13212 INV_X32 
XU53 n112 n78 NETTRAN_DUMMY_13213 NETTRAN_DUMMY_13214 CLKBUF_X1 
XU54 n80 n79 NETTRAN_DUMMY_13215 NETTRAN_DUMMY_13216 CLKBUF_X1 
XU55 n78 n80 NETTRAN_DUMMY_13217 NETTRAN_DUMMY_13218 INV_X32 
XU56 n79 p[26] NETTRAN_DUMMY_13219 NETTRAN_DUMMY_13220 INV_X32 
XU57 n111 n82 NETTRAN_DUMMY_13221 NETTRAN_DUMMY_13222 CLKBUF_X1 
XU58 n84 n83 NETTRAN_DUMMY_13223 NETTRAN_DUMMY_13224 CLKBUF_X1 
XU59 n82 n84 NETTRAN_DUMMY_13225 NETTRAN_DUMMY_13226 INV_X32 
XU60 n83 p[25] NETTRAN_DUMMY_13227 NETTRAN_DUMMY_13228 INV_X32 
XU61 n123 n86 NETTRAN_DUMMY_13229 NETTRAN_DUMMY_13230 CLKBUF_X1 
XU62 n88 n87 NETTRAN_DUMMY_13231 NETTRAN_DUMMY_13232 CLKBUF_X1 
XU63 n86 n88 NETTRAN_DUMMY_13233 NETTRAN_DUMMY_13234 INV_X32 
XU64 n87 p[24] NETTRAN_DUMMY_13235 NETTRAN_DUMMY_13236 INV_X32 
XU65 n122 n90 NETTRAN_DUMMY_13237 NETTRAN_DUMMY_13238 CLKBUF_X1 
XU66 n92 n91 NETTRAN_DUMMY_13239 NETTRAN_DUMMY_13240 CLKBUF_X1 
XU67 n90 n92 NETTRAN_DUMMY_13241 NETTRAN_DUMMY_13242 INV_X32 
XU68 n91 p[23] NETTRAN_DUMMY_13243 NETTRAN_DUMMY_13244 INV_X32 
XU69 n121 n94 NETTRAN_DUMMY_13245 NETTRAN_DUMMY_13246 CLKBUF_X1 
XU70 n96 n95 NETTRAN_DUMMY_13247 NETTRAN_DUMMY_13248 CLKBUF_X1 
XU71 n94 n96 NETTRAN_DUMMY_13249 NETTRAN_DUMMY_13250 INV_X32 
XU72 n95 p[22] NETTRAN_DUMMY_13251 NETTRAN_DUMMY_13252 INV_X32 
XU73 n101 p[21] NETTRAN_DUMMY_13253 NETTRAN_DUMMY_13254 BUF_X1 
XU74 n100 n99 NETTRAN_DUMMY_13255 NETTRAN_DUMMY_13256 CLKBUF_X1 
XU75 n120 n100 NETTRAN_DUMMY_13257 NETTRAN_DUMMY_13258 INV_X32 
XU76 n99 n101 NETTRAN_DUMMY_13259 NETTRAN_DUMMY_13260 INV_X32 
XU77 n105 p[20] NETTRAN_DUMMY_13261 NETTRAN_DUMMY_13262 BUF_X1 
XU78 n104 n103 NETTRAN_DUMMY_13263 NETTRAN_DUMMY_13264 CLKBUF_X1 
XU79 n119 n104 NETTRAN_DUMMY_13265 NETTRAN_DUMMY_13266 INV_X32 
XU80 n103 n105 NETTRAN_DUMMY_13267 NETTRAN_DUMMY_13268 INV_X32 
XU81 sum[25] n124 NETTRAN_DUMMY_13269 NETTRAN_DUMMY_13270 BUF_X1 
Xadd_69 sum[37] sum[36] sum[35] sum[34] sum[33] sum[32] sum[31] sum[30] sum[29] 
+ sum[28] sum[27] sum[26] sum[25] sum[24] sum[23] sum[22] sum[21] sum[20] sum[19] 
+ sum[18] sum[17] sum[16] sum[15] sum[14] sum[13] sum[12] sum[11] sum[10] sum[9] 
+ sum[8] sum[7] sum[6] sum[5] sum[4] sum[3] sum[2] sum[1] sum[0] VSS NETTRAN_DUMMY_13271 
+ prod[33] prod[33] prod[33] prod[33] prod[33] prod[32] prod[31] prod[30] prod[29] 
+ prod[28] prod[27] prod[26] prod[25] prod[24] prod[23] prod[22] prod[21] prod[20] 
+ prod[19] prod[18] prod[17] prod[16] prod[15] prod[14] prod[13] prod[12] prod[11] 
+ prod[10] prod[9] prod[8] prod[7] prod[6] prod[5] prod[4] prod[3] prod[2] prod[1] 
+ prod[0] c_reg[36] c_reg[36] c_reg[35] c_reg[34] c_reg[33] c_reg[32] c_reg[31] 
+ c_reg[30] c_reg[29] c_reg[28] c_reg[27] c_reg[26] c_reg[25] c_reg[24] c_reg[23] 
+ c_reg[22] c_reg[21] c_reg[20] c_reg[19] c_reg[18] c_reg[17] c_reg[16] c_reg[15] 
+ c_reg[14] c_reg[13] c_reg[12] c_reg[11] c_reg[10] c_reg[9] c_reg[8] c_reg[7] c_reg[6] 
+ c_reg[5] c_reg[4] c_reg[3] c_reg[2] c_reg[1] c_reg[0] gng_smul_16_18_sadd_37_DW01_add_0 
Xmult_66 N33 N320 N310 N301 N290 N28 N27 N26 N25 N24 N23 N22 N21 N201 N19 N18 N17 
+ N16 N15 N14 N13 N12 N11 N102 N9 N8 N7 N6 N5 N4 N300 N200 N1000 N0 VDD n302 b_reg[16] 
+ b_reg[15] b_reg[14] b_reg[13] b_reg[12] b_reg[11] b_reg[10] b_reg[9] b_reg[8] 
+ b_reg[7] b_reg[6] b_reg[5] b_reg[4] b_reg[3] b_reg[2] b_reg[1] b_reg[0] n330 a_reg[14] 
+ a_reg[13] a_reg[12] a_reg[11] a_reg[10] a_reg[9] a_reg[8] a_reg[7] a_reg[6] a_reg[5] 
+ a_reg[4] a_reg[3] a_reg[2] a_reg[1] a_reg[0] gng_smul_16_18_sadd_37_DW02_mult_0 
.ENDS

.SUBCKT gng_smul_16_18 p[33] p[32] p[31] p[30] p[29] p[28] p[27] p[26] p[25] p[24] 
+ p[23] p[22] p[21] p[20] p[19] p[18] p[17] p[16] p[15] p[14] p[13] p[12] p[11] 
+ p[10] p[9] p[8] p[7] p[6] p[5] p[4] p[3] p[2] p[1] p[0] clk b[17] b[16] b[15] 
+ b[14] b[13] b[12] b[11] b[10] b[9] b[8] b[7] b[6] b[5] b[4] b[3] b[2] b[1] b[0] 
+ a[15] a[14] a[13] a[12] a[11] a[10] a[9] a[8] a[7] a[6] a[5] a[4] a[3] a[2] a[1] 
+ a[0] 
XLOGIC0_X1_U0 LOGIC0_X1_U0_net NETTRAN_DUMMY_13272 NETTRAN_DUMMY_13273 LOGIC0_X1 
Xprod_reg_19_ N19 n1_G3B1I4 p[19] NETTRAN_DUMMY_13274 NETTRAN_DUMMY_13275 NETTRAN_DUMMY_13276 DFF_X1 
Xprod_reg_20_ N20 n1_G3B1I4 p[20] NETTRAN_DUMMY_13277 NETTRAN_DUMMY_13278 NETTRAN_DUMMY_13279 DFF_X1 
Xprod_reg_21_ N21 n1_G3B1I3 p[21] NETTRAN_DUMMY_13280 NETTRAN_DUMMY_13281 NETTRAN_DUMMY_13282 DFF_X1 
Xprod_reg_22_ N22 n1_G3B1I2 p[22] NETTRAN_DUMMY_13283 NETTRAN_DUMMY_13284 NETTRAN_DUMMY_13285 DFF_X1 
Xprod_reg_23_ N23 n1_G3B1I2 p[23] NETTRAN_DUMMY_13286 NETTRAN_DUMMY_13287 NETTRAN_DUMMY_13288 DFF_X1 
Xprod_reg_24_ N24 n1_G3B1I2 p[24] NETTRAN_DUMMY_13289 NETTRAN_DUMMY_13290 NETTRAN_DUMMY_13291 DFF_X1 
Xprod_reg_25_ N25 n1_G3B1I2 p[25] NETTRAN_DUMMY_13292 NETTRAN_DUMMY_13293 NETTRAN_DUMMY_13294 DFF_X1 
Xprod_reg_26_ N26 n1_G3B1I3 p[26] NETTRAN_DUMMY_13295 NETTRAN_DUMMY_13296 NETTRAN_DUMMY_13297 DFF_X1 
Xprod_reg_27_ N27 n1_G3B1I3 p[27] NETTRAN_DUMMY_13298 NETTRAN_DUMMY_13299 NETTRAN_DUMMY_13300 DFF_X1 
Xprod_reg_28_ N28 n1_G3B1I3 p[28] NETTRAN_DUMMY_13301 NETTRAN_DUMMY_13302 NETTRAN_DUMMY_13303 DFF_X1 
Xprod_reg_29_ N29 n1_G3B1I4 p[29] NETTRAN_DUMMY_13304 NETTRAN_DUMMY_13305 NETTRAN_DUMMY_13306 DFF_X1 
Xprod_reg_30_ N30 n1 p[30] NETTRAN_DUMMY_13307 NETTRAN_DUMMY_13308 NETTRAN_DUMMY_13309 DFF_X1 
Xprod_reg_31_ N31 n1 p[31] NETTRAN_DUMMY_13310 NETTRAN_DUMMY_13311 NETTRAN_DUMMY_13312 DFF_X1 
Xprod_reg_32_ N32 clk p[32] NETTRAN_DUMMY_13313 NETTRAN_DUMMY_13314 NETTRAN_DUMMY_13315 DFF_X1 
Xb_reg_reg_0_ b[0] clk b_reg[0] NETTRAN_DUMMY_13316 NETTRAN_DUMMY_13317 NETTRAN_DUMMY_13318 DFF_X1 
Xb_reg_reg_1_ b[1] clk b_reg[1] NETTRAN_DUMMY_13319 NETTRAN_DUMMY_13320 NETTRAN_DUMMY_13321 DFF_X1 
Xb_reg_reg_2_ b[2] n2_G3B1I1 b_reg[2] NETTRAN_DUMMY_13322 NETTRAN_DUMMY_13323 NETTRAN_DUMMY_13324 DFF_X1 
Xb_reg_reg_3_ b[3] n2_G3B1I2 b_reg[3] NETTRAN_DUMMY_13325 NETTRAN_DUMMY_13326 NETTRAN_DUMMY_13327 DFF_X1 
Xb_reg_reg_4_ b[4] n2_G3B1I4 b_reg[4] NETTRAN_DUMMY_13328 NETTRAN_DUMMY_13329 NETTRAN_DUMMY_13330 DFF_X1 
Xb_reg_reg_5_ b[5] n1_G3B1I3 b_reg[5] NETTRAN_DUMMY_13331 NETTRAN_DUMMY_13332 NETTRAN_DUMMY_13333 DFF_X1 
Xb_reg_reg_6_ b[6] n1_G3B1I3 b_reg[6] NETTRAN_DUMMY_13334 NETTRAN_DUMMY_13335 NETTRAN_DUMMY_13336 DFF_X1 
Xb_reg_reg_7_ b[7] n1_G3B1I2 b_reg[7] NETTRAN_DUMMY_13337 NETTRAN_DUMMY_13338 NETTRAN_DUMMY_13339 DFF_X1 
Xb_reg_reg_8_ b[8] n1_G3B1I3 b_reg[8] NETTRAN_DUMMY_13340 NETTRAN_DUMMY_13341 NETTRAN_DUMMY_13342 DFF_X1 
Xb_reg_reg_9_ b[9] n1_G3B1I3 b_reg[9] NETTRAN_DUMMY_13343 NETTRAN_DUMMY_13344 NETTRAN_DUMMY_13345 DFF_X1 
Xb_reg_reg_10_ b[10] n1_G3B1I3 b_reg[10] NETTRAN_DUMMY_13346 NETTRAN_DUMMY_13347 
+ NETTRAN_DUMMY_13348 DFF_X1 
Xb_reg_reg_11_ b[11] n1_G3B1I4 b_reg[11] NETTRAN_DUMMY_13349 NETTRAN_DUMMY_13350 
+ NETTRAN_DUMMY_13351 DFF_X1 
Xb_reg_reg_12_ b[12] n1_G3B1I4 b_reg[12] NETTRAN_DUMMY_13352 NETTRAN_DUMMY_13353 
+ NETTRAN_DUMMY_13354 DFF_X1 
Xb_reg_reg_13_ b[13] n1_G3B1I4 b_reg[13] NETTRAN_DUMMY_13355 NETTRAN_DUMMY_13356 
+ NETTRAN_DUMMY_13357 DFF_X1 
Xb_reg_reg_14_ b[14] n1 b_reg[14] NETTRAN_DUMMY_13358 NETTRAN_DUMMY_13359 NETTRAN_DUMMY_13360 DFF_X1 
Xb_reg_reg_15_ b[15] n1 b_reg[15] NETTRAN_DUMMY_13361 NETTRAN_DUMMY_13362 NETTRAN_DUMMY_13363 DFF_X1 
Xb_reg_reg_16_ b[16] n1 b_reg[16] NETTRAN_DUMMY_13364 NETTRAN_DUMMY_13365 NETTRAN_DUMMY_13366 DFF_X1 
Xb_reg_reg_17_ b[17] n2_G3B1I4 b_reg[17] NETTRAN_DUMMY_13367 NETTRAN_DUMMY_13368 
+ NETTRAN_DUMMY_13369 DFF_X1 
Xa_reg_reg_0_ a[0] n2_G3B1I2 a_reg[0] NETTRAN_DUMMY_13370 NETTRAN_DUMMY_13371 NETTRAN_DUMMY_13372 DFF_X1 
Xa_reg_reg_1_ a[1] n2_G3B1I1 a_reg[1] NETTRAN_DUMMY_13373 NETTRAN_DUMMY_13374 NETTRAN_DUMMY_13375 DFF_X1 
Xa_reg_reg_2_ a[2] n2_G3B1I2 a_reg[2] NETTRAN_DUMMY_13376 NETTRAN_DUMMY_13377 NETTRAN_DUMMY_13378 DFF_X1 
Xa_reg_reg_3_ a[3] n2_G3B1I2 a_reg[3] NETTRAN_DUMMY_13379 NETTRAN_DUMMY_13380 NETTRAN_DUMMY_13381 DFF_X1 
Xa_reg_reg_4_ a[4] n2_G3B1I2 a_reg[4] NETTRAN_DUMMY_13382 NETTRAN_DUMMY_13383 NETTRAN_DUMMY_13384 DFF_X1 
Xa_reg_reg_5_ a[5] n2_G3B1I1 a_reg[5] NETTRAN_DUMMY_13385 NETTRAN_DUMMY_13386 NETTRAN_DUMMY_13387 DFF_X1 
Xa_reg_reg_6_ a[6] n2_G3B1I4 a_reg[6] NETTRAN_DUMMY_13388 NETTRAN_DUMMY_13389 NETTRAN_DUMMY_13390 DFF_X1 
Xa_reg_reg_7_ a[7] n2_G3B1I4 a_reg[7] NETTRAN_DUMMY_13391 NETTRAN_DUMMY_13392 NETTRAN_DUMMY_13393 DFF_X1 
Xa_reg_reg_8_ a[8] n2_G3B1I4 a_reg[8] NETTRAN_DUMMY_13394 NETTRAN_DUMMY_13395 NETTRAN_DUMMY_13396 DFF_X1 
Xa_reg_reg_9_ a[9] n1 a_reg[9] NETTRAN_DUMMY_13397 NETTRAN_DUMMY_13398 NETTRAN_DUMMY_13399 DFF_X1 
Xa_reg_reg_10_ a[10] n2_G3B1I1 a_reg[10] NETTRAN_DUMMY_13400 NETTRAN_DUMMY_13401 
+ NETTRAN_DUMMY_13402 DFF_X1 
Xa_reg_reg_11_ a[11] n2_G3B1I1 a_reg[11] NETTRAN_DUMMY_13403 NETTRAN_DUMMY_13404 
+ NETTRAN_DUMMY_13405 DFF_X1 
Xa_reg_reg_12_ a[12] n2_G3B1I4 a_reg[12] NETTRAN_DUMMY_13406 NETTRAN_DUMMY_13407 
+ NETTRAN_DUMMY_13408 DFF_X1 
Xa_reg_reg_13_ a[13] n2_G3B1I4 a_reg[13] NETTRAN_DUMMY_13409 NETTRAN_DUMMY_13410 
+ NETTRAN_DUMMY_13411 DFF_X1 
Xa_reg_reg_14_ a[14] n2_G3B1I4 a_reg[14] NETTRAN_DUMMY_13412 NETTRAN_DUMMY_13413 
+ NETTRAN_DUMMY_13414 DFF_X1 
Xa_reg_reg_15_ LOGIC0_X1_U0_net n2_G3B1I2 a_reg[15] NETTRAN_DUMMY_13415 NETTRAN_DUMMY_13416 
+ NETTRAN_DUMMY_13417 DFF_X1 
XU1 clk n1 NETTRAN_DUMMY_13418 NETTRAN_DUMMY_13419 BUF_X32 
XCLKBUF_X1_G3B1I21 n1 n1_G3B1I2 NETTRAN_DUMMY_13420 NETTRAN_DUMMY_13421 CLKBUF_X1 
XCLKBUF_X1_G3B1I4 clk n2_G3B1I4 NETTRAN_DUMMY_13422 NETTRAN_DUMMY_13423 CLKBUF_X2 
XCLKBUF_X1_G3B1I31 n1 n1_G3B1I3 NETTRAN_DUMMY_13424 NETTRAN_DUMMY_13425 CLKBUF_X2 
XCLKBUF_X1_G3B1I41 n1 n1_G3B1I4 NETTRAN_DUMMY_13426 NETTRAN_DUMMY_13427 CLKBUF_X2 
XCLKBUF_X1_G3B1I1 clk n2_G3B1I1 NETTRAN_DUMMY_13428 NETTRAN_DUMMY_13429 CLKBUF_X2 
XCLKBUF_X1_G3B1I2 clk n2_G3B1I2 NETTRAN_DUMMY_13430 NETTRAN_DUMMY_13431 CLKBUF_X2 
Xmult_60 N33 N32 N31 N30 N29 N28 N27 N26 N25 N24 N23 N22 N21 N20 N19 N18 N17 N16 
+ N15 N14 N13 N12 N11 N101 N9 N8 N7 N6 N5 N4 N3 N2 N100 N0 VDD b_reg[17] b_reg[16] 
+ b_reg[15] b_reg[14] b_reg[13] b_reg[12] b_reg[11] b_reg[10] b_reg[9] b_reg[8] 
+ b_reg[7] b_reg[6] b_reg[5] b_reg[4] b_reg[3] b_reg[2] b_reg[1] b_reg[0] a_reg[15] 
+ a_reg[14] a_reg[13] a_reg[12] a_reg[11] a_reg[10] a_reg[9] a_reg[8] a_reg[7] a_reg[6] 
+ a_reg[5] a_reg[4] a_reg[3] a_reg[2] a_reg[1] a_reg[0] gng_smul_16_18_DW02_mult_0 
.ENDS

.SUBCKT gng_interp clk rstn valid_in valid_out IN0 IN1 data_out[15] data_out[14] 
+ data_out[13] data_out[12] data_out[11] data_out[10] data_out[9] data_out[8] data_out[7] 
+ data_out[6] data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] 
+ data_in[63] data_in[62] data_in[61] data_in[60] data_in[59] data_in[58] data_in[57] 
+ data_in[56] data_in[55] data_in[54] data_in[53] data_in[52] data_in[51] data_in[50] 
+ data_in[49] data_in[48] data_in[47] data_in[46] data_in[45] data_in[44] data_in[43] 
+ data_in[42] data_in[41] data_in[40] data_in[39] data_in[38] data_in[37] data_in[36] 
+ data_in[35] data_in[34] data_in[33] data_in[32] data_in[31] data_in[30] data_in[29] 
+ data_in[28] data_in[27] data_in[26] data_in[25] data_in[24] data_in[23] data_in[22] 
+ data_in[21] data_in[20] data_in[19] data_in[18] data_in[17] data_in[16] data_in[15] 
+ data_in[14] data_in[13] data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] 
+ data_in[7] data_in[6] data_in[5] data_in[4] data_in[3] data_in[2] data_in[1] data_in[0] 
+ IN2 clk_cts_3 
XU153 n132 n7310 NETTRAN_DUMMY_13432 NETTRAN_DUMMY_13433 CLKBUF_X2 
XU152 n204 n7210 NETTRAN_DUMMY_13434 NETTRAN_DUMMY_13435 BUF_X1 
XU150 n142 n7011 NETTRAN_DUMMY_13436 NETTRAN_DUMMY_13437 BUF_X2 
XU148 n208 n6810 NETTRAN_DUMMY_13438 NETTRAN_DUMMY_13439 BUF_X2 
Xx_r2_reg_7_ n1303 n10_G2B1I4 x_r2[7] NETTRAN_DUMMY_13440 NETTRAN_DUMMY_13441 NETTRAN_DUMMY_13442 DFF_X1 
Xx_r1_reg_7_ n201 n6_G2B1I4 x_r1[7] NETTRAN_DUMMY_13443 NETTRAN_DUMMY_13444 NETTRAN_DUMMY_13445 DFF_X1 
Xx_r3_reg_8_ n1293 n10_G2B1I3 x_r3[8] NETTRAN_DUMMY_13446 NETTRAN_DUMMY_13447 NETTRAN_DUMMY_13448 DFF_X1 
Xx_r2_reg_8_ n209 n10_G2B1I4 x_r2[8] NETTRAN_DUMMY_13449 NETTRAN_DUMMY_13450 NETTRAN_DUMMY_13451 DFF_X1 
Xx_r1_reg_8_ n1334 n60 x_r1[8] NETTRAN_DUMMY_13452 NETTRAN_DUMMY_13453 NETTRAN_DUMMY_13454 DFF_X1 
Xx_r3_reg_9_ n1280 n8_G2B1I2 x_r3[9] NETTRAN_DUMMY_13455 NETTRAN_DUMMY_13456 NETTRAN_DUMMY_13457 DFF_X1 
Xx_r2_reg_9_ n1276 n8_G2B1I7 x_r2[9] NETTRAN_DUMMY_13458 NETTRAN_DUMMY_13459 NETTRAN_DUMMY_13460 DFF_X1 
Xx_r1_reg_9_ n1307 n8_G2B1I2 x_r1[9] NETTRAN_DUMMY_13461 NETTRAN_DUMMY_13462 NETTRAN_DUMMY_13463 DFF_X1 
Xx_r3_reg_10_ n1266 n10_G2B1I4 x_r3[10] NETTRAN_DUMMY_13464 NETTRAN_DUMMY_13465 
+ NETTRAN_DUMMY_13466 DFF_X1 
Xx_r2_reg_10_ n1262 n6_G2B1I5 x_r2[10] NETTRAN_DUMMY_13467 NETTRAN_DUMMY_13468 NETTRAN_DUMMY_13469 DFF_X1 
Xx_r1_reg_10_ n200 n6_G2B1I4 x_r1[10] NETTRAN_DUMMY_13470 NETTRAN_DUMMY_13471 NETTRAN_DUMMY_13472 DFF_X1 
Xx_r3_reg_11_ n1253 n10_G2B1I4 x_r3[11] NETTRAN_DUMMY_13473 NETTRAN_DUMMY_13474 
+ NETTRAN_DUMMY_13475 DFF_X1 
Xx_r2_reg_11_ n1249 n6_G2B1I5 x_r2[11] NETTRAN_DUMMY_13476 NETTRAN_DUMMY_13477 NETTRAN_DUMMY_13478 DFF_X1 
Xx_r1_reg_11_ n198 n6_G2B1I4 x_r1[11] NETTRAN_DUMMY_13479 NETTRAN_DUMMY_13480 NETTRAN_DUMMY_13481 DFF_X1 
Xx_r3_reg_12_ n1239 n10_G2B1I2 x_r3[12] NETTRAN_DUMMY_13482 NETTRAN_DUMMY_13483 
+ NETTRAN_DUMMY_13484 DFF_X1 
Xx_r2_reg_12_ n1235 n10_G2B1I4 x_r2[12] NETTRAN_DUMMY_13485 NETTRAN_DUMMY_13486 
+ NETTRAN_DUMMY_13487 DFF_X1 
Xx_r1_reg_12_ n1970 n6_G2B1I4 x_r1[12] NETTRAN_DUMMY_13488 NETTRAN_DUMMY_13489 NETTRAN_DUMMY_13490 DFF_X1 
Xx_r3_reg_13_ n1226 n10_G2B1I3 x_r3[13] NETTRAN_DUMMY_13491 NETTRAN_DUMMY_13492 
+ NETTRAN_DUMMY_13493 DFF_X1 
Xx_r2_reg_13_ n1222 n10_G2B1I2 x_r2[13] NETTRAN_DUMMY_13494 NETTRAN_DUMMY_13495 
+ NETTRAN_DUMMY_13496 DFF_X1 
Xx_r1_reg_13_ n1950 n6_G2B1I3 x_r1[13] NETTRAN_DUMMY_13497 NETTRAN_DUMMY_13498 NETTRAN_DUMMY_13499 DFF_X1 
Xx_r3_reg_14_ n1212 n10_G2B1I2 x_r3[14] NETTRAN_DUMMY_13500 NETTRAN_DUMMY_13501 
+ NETTRAN_DUMMY_13502 DFF_X1 
Xx_r2_reg_14_ n1208 n10_G2B1I2 x_r2[14] NETTRAN_DUMMY_13503 NETTRAN_DUMMY_13504 
+ NETTRAN_DUMMY_13505 DFF_X1 
Xx_r1_reg_14_ n1940 n6_G2B1I3 x_r1[14] NETTRAN_DUMMY_13506 NETTRAN_DUMMY_13507 NETTRAN_DUMMY_13508 DFF_X1 
Xx_reg_0_ n1195 n11_G2B1I7 NETTRAN_DUMMY_13509 n59 NETTRAN_DUMMY_13510 NETTRAN_DUMMY_13511 DFF_X1 
Xx_reg_1_ n1191 n11_G2B1I7 NETTRAN_DUMMY_13512 n6110 NETTRAN_DUMMY_13513 NETTRAN_DUMMY_13514 DFF_X1 
Xx_reg_2_ n1190 n11_G2B1I6 NETTRAN_DUMMY_13515 n630 NETTRAN_DUMMY_13516 NETTRAN_DUMMY_13517 DFF_X1 
Xx_reg_3_ N80 n11_G2B1I6 NETTRAN_DUMMY_13518 n650 NETTRAN_DUMMY_13519 NETTRAN_DUMMY_13520 DFF_X1 
Xx_reg_4_ n1186 n11_G2B1I1 NETTRAN_DUMMY_13521 n670 NETTRAN_DUMMY_13522 NETTRAN_DUMMY_13523 DFF_X1 
Xx_reg_5_ n1182 n11_G2B1I4 NETTRAN_DUMMY_13524 n690 NETTRAN_DUMMY_13525 NETTRAN_DUMMY_13526 DFF_X1 
Xx_reg_6_ n1178 n11_G2B1I5 NETTRAN_DUMMY_13527 n711 NETTRAN_DUMMY_13528 NETTRAN_DUMMY_13529 DFF_X1 
Xx_reg_7_ n1174 n11_G2B1I3 NETTRAN_DUMMY_13530 n730 NETTRAN_DUMMY_13531 NETTRAN_DUMMY_13532 DFF_X1 
Xx_reg_8_ n1167 n11_G2B1I6 NETTRAN_DUMMY_13533 n750 NETTRAN_DUMMY_13534 NETTRAN_DUMMY_13535 DFF_X1 
Xx_reg_9_ n1166 n2 NETTRAN_DUMMY_13536 n770 NETTRAN_DUMMY_13537 NETTRAN_DUMMY_13538 DFF_X1 
Xx_reg_10_ n1163 n11_G2B1I2 NETTRAN_DUMMY_13539 n790 NETTRAN_DUMMY_13540 NETTRAN_DUMMY_13541 DFF_X1 
Xx_reg_11_ n1159 n11_G2B1I3 NETTRAN_DUMMY_13542 n811 NETTRAN_DUMMY_13543 NETTRAN_DUMMY_13544 DFF_X1 
Xx_reg_12_ n1157 n11_G2B1I3 NETTRAN_DUMMY_13545 n830 NETTRAN_DUMMY_13546 NETTRAN_DUMMY_13547 DFF_X1 
Xx_reg_13_ n1153 n11_G2B1I3 NETTRAN_DUMMY_13548 n850 NETTRAN_DUMMY_13549 NETTRAN_DUMMY_13550 DFF_X1 
Xx_reg_14_ n1149 n11_G2B1I3 NETTRAN_DUMMY_13551 n870 NETTRAN_DUMMY_13552 NETTRAN_DUMMY_13553 DFF_X1 
Xoffset_reg_0_ n1142 n6 offset[0] NETTRAN_DUMMY_13554 NETTRAN_DUMMY_13555 NETTRAN_DUMMY_13556 DFF_X1 
Xoffset_reg_1_ n1141 n8_G2B1I7 offset[1] NETTRAN_DUMMY_13557 NETTRAN_DUMMY_13558 
+ NETTRAN_DUMMY_13559 DFF_X1 
Xmask_reg_0_ n1134 n11_G2B1I7 NETTRAN_DUMMY_13560 n6000 NETTRAN_DUMMY_13561 NETTRAN_DUMMY_13562 DFF_X1 
Xmask_reg_1_ n1129 n11_G2B1I7 NETTRAN_DUMMY_13563 n6200 NETTRAN_DUMMY_13564 NETTRAN_DUMMY_13565 DFF_X1 
Xmask_reg_2_ N620 n11_G2B1I5 NETTRAN_DUMMY_13566 n640 NETTRAN_DUMMY_13567 NETTRAN_DUMMY_13568 DFF_X1 
Xmask_reg_3_ N63 n11_G2B1I6 NETTRAN_DUMMY_13569 n660 NETTRAN_DUMMY_13570 NETTRAN_DUMMY_13571 DFF_X1 
Xmask_reg_4_ n1109 n11_G2B1I6 NETTRAN_DUMMY_13572 n680 NETTRAN_DUMMY_13573 NETTRAN_DUMMY_13574 DFF_X1 
Xmask_reg_5_ n1103 n11_G2B1I5 NETTRAN_DUMMY_13575 n7000 NETTRAN_DUMMY_13576 NETTRAN_DUMMY_13577 DFF_X1 
Xmask_reg_6_ N66 n11_G2B1I5 NETTRAN_DUMMY_13578 n720 NETTRAN_DUMMY_13579 NETTRAN_DUMMY_13580 DFF_X1 
Xmask_reg_7_ N67 n11_G2B1I2 NETTRAN_DUMMY_13581 n740 NETTRAN_DUMMY_13582 NETTRAN_DUMMY_13583 DFF_X1 
Xmask_reg_8_ N68 n11_G2B1I6 NETTRAN_DUMMY_13584 n760 NETTRAN_DUMMY_13585 NETTRAN_DUMMY_13586 DFF_X1 
Xmask_reg_9_ N69 n11_G2B1I4 NETTRAN_DUMMY_13587 n780 NETTRAN_DUMMY_13588 NETTRAN_DUMMY_13589 DFF_X1 
Xmask_reg_10_ n1085 n6_G2B1I3 NETTRAN_DUMMY_13590 n800 NETTRAN_DUMMY_13591 NETTRAN_DUMMY_13592 DFF_X1 
Xmask_reg_11_ N71 n11_G2B1I2 NETTRAN_DUMMY_13593 n820 NETTRAN_DUMMY_13594 NETTRAN_DUMMY_13595 DFF_X1 
Xmask_reg_12_ N72 n11_G2B1I5 NETTRAN_DUMMY_13596 n840 NETTRAN_DUMMY_13597 NETTRAN_DUMMY_13598 DFF_X1 
Xmask_reg_13_ N73 n11_G2B1I2 NETTRAN_DUMMY_13599 n860 NETTRAN_DUMMY_13600 NETTRAN_DUMMY_13601 DFF_X1 
Xmask_reg_14_ n1083 n11_G2B1I2 NETTRAN_DUMMY_13602 n880 NETTRAN_DUMMY_13603 NETTRAN_DUMMY_13604 DFF_X1 
Xnum_lzd_r_reg_0_ n1920 n11_G2B1I4 num_lzd_r[0] n1110 NETTRAN_DUMMY_13605 NETTRAN_DUMMY_13606 DFF_X2 
Xnum_lzd_r_reg_1_ n1082 n11_G2B1I4 num_lzd_r[1] n1010 NETTRAN_DUMMY_13607 NETTRAN_DUMMY_13608 DFF_X1 
Xnum_lzd_r_reg_2_ n1081 n11_G2B1I4 num_lzd_r[2] n910 NETTRAN_DUMMY_13609 NETTRAN_DUMMY_13610 DFF_X1 
Xnum_lzd_r_reg_3_ n1079 n11_G2B1I3 num_lzd_r[3] n810 NETTRAN_DUMMY_13611 NETTRAN_DUMMY_13612 DFF_X1 
Xnum_lzd_r_reg_4_ n1075 n11_G2B1I4 num_lzd_r[4] n710 NETTRAN_DUMMY_13613 NETTRAN_DUMMY_13614 DFF_X1 
Xnum_lzd_r_reg_5_ n1073 n11_G2B1I4 num_lzd_r[5] NETTRAN_DUMMY_13615 NETTRAN_DUMMY_13616 
+ NETTRAN_DUMMY_13617 DFF_X1 
Xc0_r2_reg_8_ n1071 n7_G2B1I1 c0_r2[8] NETTRAN_DUMMY_13618 NETTRAN_DUMMY_13619 NETTRAN_DUMMY_13620 DFF_X1 
Xc0_r1_reg_8_ c0[8] n7_G2B1I1 c0_r1[8] NETTRAN_DUMMY_13621 NETTRAN_DUMMY_13622 NETTRAN_DUMMY_13623 DFF_X1 
Xc0_r4_reg_9_ n1066 n7_G2B1I4 c0_r4[9] NETTRAN_DUMMY_13624 NETTRAN_DUMMY_13625 NETTRAN_DUMMY_13626 DFF_X1 
Xc0_r3_reg_9_ n1062 n7_G2B1I4 c0_r3[9] NETTRAN_DUMMY_13627 NETTRAN_DUMMY_13628 NETTRAN_DUMMY_13629 DFF_X1 
Xc0_r2_reg_9_ n1880 n7_G2B1I4 c0_r2[9] NETTRAN_DUMMY_13630 NETTRAN_DUMMY_13631 NETTRAN_DUMMY_13632 DFF_X1 
Xc0_r1_reg_9_ c0[9] n62 c0_r1[9] NETTRAN_DUMMY_13633 NETTRAN_DUMMY_13634 NETTRAN_DUMMY_13635 DFF_X1 
Xc0_r4_reg_10_ n1049 n62 c0_r4[10] NETTRAN_DUMMY_13636 NETTRAN_DUMMY_13637 NETTRAN_DUMMY_13638 DFF_X1 
Xc0_r3_reg_10_ n1048 n62_G2B1I2 c0_r3[10] NETTRAN_DUMMY_13639 NETTRAN_DUMMY_13640 
+ NETTRAN_DUMMY_13641 DFF_X1 
Xc0_r2_reg_10_ n1044 n62_G2B1I2 c0_r2[10] NETTRAN_DUMMY_13642 NETTRAN_DUMMY_13643 
+ NETTRAN_DUMMY_13644 DFF_X1 
Xc0_r1_reg_10_ c0[10] n63_G2B1I2 c0_r1[10] NETTRAN_DUMMY_13645 NETTRAN_DUMMY_13646 
+ NETTRAN_DUMMY_13647 DFF_X1 
Xc0_r4_reg_11_ n1039 n6_G2B1I5 c0_r4[11] NETTRAN_DUMMY_13648 NETTRAN_DUMMY_13649 
+ NETTRAN_DUMMY_13650 DFF_X1 
Xc0_r3_reg_11_ n1035 n6_G2B1I5 c0_r3[11] NETTRAN_DUMMY_13651 NETTRAN_DUMMY_13652 
+ NETTRAN_DUMMY_13653 DFF_X1 
Xc0_r2_reg_11_ n1031 n6_G2B1I3 c0_r2[11] NETTRAN_DUMMY_13654 NETTRAN_DUMMY_13655 
+ NETTRAN_DUMMY_13656 DFF_X1 
Xc0_r1_reg_11_ c0[11] n6_G2B1I3 c0_r1[11] NETTRAN_DUMMY_13657 NETTRAN_DUMMY_13658 
+ NETTRAN_DUMMY_13659 DFF_X1 
Xc0_r4_reg_12_ n1026 n6_G2B1I5 c0_r4[12] NETTRAN_DUMMY_13660 NETTRAN_DUMMY_13661 
+ NETTRAN_DUMMY_13662 DFF_X1 
Xc0_r3_reg_12_ n1022 n6_G2B1I3 c0_r3[12] NETTRAN_DUMMY_13663 NETTRAN_DUMMY_13664 
+ NETTRAN_DUMMY_13665 DFF_X1 
Xc0_r2_reg_12_ n1870 n6_G2B1I3 c0_r2[12] NETTRAN_DUMMY_13666 NETTRAN_DUMMY_13667 
+ NETTRAN_DUMMY_13668 DFF_X1 
Xc0_r1_reg_12_ c0[12] n6 c0_r1[12] NETTRAN_DUMMY_13669 NETTRAN_DUMMY_13670 NETTRAN_DUMMY_13671 DFF_X1 
Xc0_r4_reg_13_ n1013 n60_G2B1I5 c0_r4[13] NETTRAN_DUMMY_13672 NETTRAN_DUMMY_13673 
+ NETTRAN_DUMMY_13674 DFF_X1 
Xc0_r3_reg_13_ n1007 n60_G2B1I5 c0_r3[13] NETTRAN_DUMMY_13675 NETTRAN_DUMMY_13676 
+ NETTRAN_DUMMY_13677 DFF_X1 
Xc0_r2_reg_13_ n1003 n60_G2B1I5 c0_r2[13] NETTRAN_DUMMY_13678 NETTRAN_DUMMY_13679 
+ NETTRAN_DUMMY_13680 DFF_X1 
Xc0_r1_reg_13_ c0[13] n11_G2B1I6 c0_r1[13] NETTRAN_DUMMY_13681 NETTRAN_DUMMY_13682 
+ NETTRAN_DUMMY_13683 DFF_X1 
Xc0_r4_reg_14_ n998 n8_G2B1I2 c0_r4[14] NETTRAN_DUMMY_13684 NETTRAN_DUMMY_13685 
+ NETTRAN_DUMMY_13686 DFF_X1 
Xc0_r3_reg_14_ n994 n8_G2B1I7 c0_r3[14] NETTRAN_DUMMY_13687 NETTRAN_DUMMY_13688 
+ NETTRAN_DUMMY_13689 DFF_X1 
Xc0_r2_reg_14_ n989 n8_G2B1I7 c0_r2[14] NETTRAN_DUMMY_13690 NETTRAN_DUMMY_13691 
+ NETTRAN_DUMMY_13692 DFF_X1 
Xc0_r1_reg_14_ c0[14] n8_G2B1I7 c0_r1[14] NETTRAN_DUMMY_13693 NETTRAN_DUMMY_13694 
+ NETTRAN_DUMMY_13695 DFF_X1 
Xc0_r4_reg_15_ n985 n11_G2B1I1 c0_r4[15] NETTRAN_DUMMY_13696 NETTRAN_DUMMY_13697 
+ NETTRAN_DUMMY_13698 DFF_X1 
Xc0_r3_reg_15_ n981 n60_G2B1I1 c0_r3[15] NETTRAN_DUMMY_13699 NETTRAN_DUMMY_13700 
+ NETTRAN_DUMMY_13701 DFF_X1 
Xc0_r2_reg_15_ n976 n60_G2B1I1 c0_r2[15] NETTRAN_DUMMY_13702 NETTRAN_DUMMY_13703 
+ NETTRAN_DUMMY_13704 DFF_X1 
Xc0_r1_reg_15_ c0[15] n60_G2B1I5 c0_r1[15] NETTRAN_DUMMY_13705 NETTRAN_DUMMY_13706 
+ NETTRAN_DUMMY_13707 DFF_X1 
Xc0_r4_reg_16_ n972 n8_G2B1I7 c0_r4[16] NETTRAN_DUMMY_13708 NETTRAN_DUMMY_13709 
+ NETTRAN_DUMMY_13710 DFF_X1 
Xc0_r3_reg_16_ n968 n8_G2B1I1 c0_r3[16] NETTRAN_DUMMY_13711 NETTRAN_DUMMY_13712 
+ NETTRAN_DUMMY_13713 DFF_X1 
Xc0_r2_reg_16_ n964 n8_G2B1I1 c0_r2[16] NETTRAN_DUMMY_13714 NETTRAN_DUMMY_13715 
+ NETTRAN_DUMMY_13716 DFF_X1 
Xc0_r1_reg_16_ c0[16] n8_G2B1I1 c0_r1[16] NETTRAN_DUMMY_13717 NETTRAN_DUMMY_13718 
+ NETTRAN_DUMMY_13719 DFF_X1 
Xc0_r4_reg_17_ n960 n11_G2B1I1 c0_r4[17] NETTRAN_DUMMY_13720 NETTRAN_DUMMY_13721 
+ NETTRAN_DUMMY_13722 DFF_X1 
Xc0_r3_reg_17_ n956 n11_G2B1I1 c0_r3[17] NETTRAN_DUMMY_13723 NETTRAN_DUMMY_13724 
+ NETTRAN_DUMMY_13725 DFF_X1 
Xc0_r2_reg_17_ n952 n11_G2B1I1 c0_r2[17] NETTRAN_DUMMY_13726 NETTRAN_DUMMY_13727 
+ NETTRAN_DUMMY_13728 DFF_X1 
Xc0_r1_reg_17_ c0[17] n11_G2B1I6 c0_r1[17] NETTRAN_DUMMY_13729 NETTRAN_DUMMY_13730 
+ NETTRAN_DUMMY_13731 DFF_X1 
Xc1_r1_reg_0_ c1[0] n11_G2B1I5 c1_r1[0] NETTRAN_DUMMY_13732 NETTRAN_DUMMY_13733 
+ NETTRAN_DUMMY_13734 DFF_X1 
Xc1_r1_reg_1_ c1[1] n6_G2B1I3 c1_r1[1] NETTRAN_DUMMY_13735 NETTRAN_DUMMY_13736 NETTRAN_DUMMY_13737 DFF_X1 
Xc1_r1_reg_2_ c1[2] n6 c1_r1[2] NETTRAN_DUMMY_13738 NETTRAN_DUMMY_13739 NETTRAN_DUMMY_13740 DFF_X1 
Xc1_r1_reg_3_ c1[3] n6_G2B1I3 c1_r1[3] NETTRAN_DUMMY_13741 NETTRAN_DUMMY_13742 NETTRAN_DUMMY_13743 DFF_X1 
Xc1_r1_reg_4_ c1[4] n6_G2B1I5 c1_r1[4] NETTRAN_DUMMY_13744 NETTRAN_DUMMY_13745 NETTRAN_DUMMY_13746 DFF_X1 
Xc1_r1_reg_5_ c1[5] n62_G2B1I2 c1_r1[5] NETTRAN_DUMMY_13747 NETTRAN_DUMMY_13748 
+ NETTRAN_DUMMY_13749 DFF_X1 
Xc1_r1_reg_6_ c1[6] n62_G2B1I2 c1_r1[6] NETTRAN_DUMMY_13750 NETTRAN_DUMMY_13751 
+ NETTRAN_DUMMY_13752 DFF_X1 
Xc1_r1_reg_7_ c1[7] n62 c1_r1[7] NETTRAN_DUMMY_13753 NETTRAN_DUMMY_13754 NETTRAN_DUMMY_13755 DFF_X1 
Xc1_r1_reg_8_ c1[8] n7_G2B1I4 c1_r1[8] NETTRAN_DUMMY_13756 NETTRAN_DUMMY_13757 NETTRAN_DUMMY_13758 DFF_X1 
Xc1_r1_reg_9_ c1[9] n7_G2B1I4 c1_r1[9] NETTRAN_DUMMY_13759 NETTRAN_DUMMY_13760 NETTRAN_DUMMY_13761 DFF_X1 
Xc1_r1_reg_10_ c1[10] n7_G2B1I4 c1_r1[10] NETTRAN_DUMMY_13762 NETTRAN_DUMMY_13763 
+ NETTRAN_DUMMY_13764 DFF_X1 
Xc1_r1_reg_11_ c1[11] n62 c1_r1[11] NETTRAN_DUMMY_13765 NETTRAN_DUMMY_13766 NETTRAN_DUMMY_13767 DFF_X1 
Xc1_r1_reg_12_ c1[12] n62_G2B1I2 c1_r1[12] NETTRAN_DUMMY_13768 NETTRAN_DUMMY_13769 
+ NETTRAN_DUMMY_13770 DFF_X1 
Xc1_r1_reg_13_ c1[13] n62_G2B1I2 c1_r1[13] NETTRAN_DUMMY_13771 NETTRAN_DUMMY_13772 
+ NETTRAN_DUMMY_13773 DFF_X1 
Xc1_r1_reg_14_ c1[14] n63_G2B1I8 c1_r1[14] NETTRAN_DUMMY_13774 NETTRAN_DUMMY_13775 
+ NETTRAN_DUMMY_13776 DFF_X1 
Xc1_r1_reg_15_ c1[15] n63_G2B1I8 c1_r1[15] NETTRAN_DUMMY_13777 NETTRAN_DUMMY_13778 
+ NETTRAN_DUMMY_13779 DFF_X1 
Xc1_r1_reg_16_ c1[16] n63_G2B1I8 c1_r1[16] NETTRAN_DUMMY_13780 NETTRAN_DUMMY_13781 
+ NETTRAN_DUMMY_13782 DFF_X1 
Xc1_r1_reg_17_ c1[17] n63_G2B1I8 c1_r1[17] NETTRAN_DUMMY_13783 NETTRAN_DUMMY_13784 
+ NETTRAN_DUMMY_13785 DFF_X1 
Xx_r4_reg_0_ n947 n6_G2B1I2 x_r4[0] NETTRAN_DUMMY_13786 NETTRAN_DUMMY_13787 NETTRAN_DUMMY_13788 DFF_X1 
Xx_r4_reg_1_ n943 n6_G2B1I2 x_r4[1] NETTRAN_DUMMY_13789 NETTRAN_DUMMY_13790 NETTRAN_DUMMY_13791 DFF_X1 
Xx_r4_reg_2_ n938 n10_G2B1I3 x_r4[2] NETTRAN_DUMMY_13792 NETTRAN_DUMMY_13793 NETTRAN_DUMMY_13794 DFF_X1 
Xx_r4_reg_3_ n934 n6_G2B1I2 x_r4[3] NETTRAN_DUMMY_13795 NETTRAN_DUMMY_13796 NETTRAN_DUMMY_13797 DFF_X1 
Xx_r4_reg_4_ n1860 n61_G2B1I1 x_r4[4] NETTRAN_DUMMY_13798 NETTRAN_DUMMY_13799 NETTRAN_DUMMY_13800 DFF_X1 
Xx_r4_reg_5_ n925 n6_G2B1I2 x_r4[5] NETTRAN_DUMMY_13801 NETTRAN_DUMMY_13802 NETTRAN_DUMMY_13803 DFF_X1 
Xx_r4_reg_6_ n1850 n61_G2B1I1 x_r4[6] NETTRAN_DUMMY_13804 NETTRAN_DUMMY_13805 NETTRAN_DUMMY_13806 DFF_X1 
Xx_r4_reg_7_ n916 n61_G2B1I1 x_r4[7] NETTRAN_DUMMY_13807 NETTRAN_DUMMY_13808 NETTRAN_DUMMY_13809 DFF_X1 
Xx_r4_reg_8_ n912 n61_G2B1I1 x_r4[8] NETTRAN_DUMMY_13810 NETTRAN_DUMMY_13811 NETTRAN_DUMMY_13812 DFF_X1 
Xx_r4_reg_9_ n906 n8_G2B1I2 x_r4[9] NETTRAN_DUMMY_13813 NETTRAN_DUMMY_13814 NETTRAN_DUMMY_13815 DFF_X1 
Xx_r4_reg_10_ n902 n10_G2B1I2 x_r4[10] NETTRAN_DUMMY_13816 NETTRAN_DUMMY_13817 NETTRAN_DUMMY_13818 DFF_X1 
Xx_r4_reg_11_ n897 n10_G2B1I2 x_r4[11] NETTRAN_DUMMY_13819 NETTRAN_DUMMY_13820 NETTRAN_DUMMY_13821 DFF_X1 
Xx_r4_reg_12_ n893 n10_G2B1I3 x_r4[12] NETTRAN_DUMMY_13822 NETTRAN_DUMMY_13823 NETTRAN_DUMMY_13824 DFF_X1 
Xx_r4_reg_13_ n888 n10_G2B1I3 x_r4[13] NETTRAN_DUMMY_13825 NETTRAN_DUMMY_13826 NETTRAN_DUMMY_13827 DFF_X1 
Xx_r4_reg_14_ n884 n10_G2B1I3 x_r4[14] NETTRAN_DUMMY_13828 NETTRAN_DUMMY_13829 NETTRAN_DUMMY_13830 DFF_X1 
Xx_r3_reg_0_ n879 n6_G2B1I2 x_r3[0] NETTRAN_DUMMY_13831 NETTRAN_DUMMY_13832 NETTRAN_DUMMY_13833 DFF_X1 
Xx_r2_reg_0_ n875 n6_G2B1I4 x_r2[0] NETTRAN_DUMMY_13834 NETTRAN_DUMMY_13835 NETTRAN_DUMMY_13836 DFF_X1 
Xx_r1_reg_0_ n141 n11_G2B1I5 x_r1[0] NETTRAN_DUMMY_13837 NETTRAN_DUMMY_13838 NETTRAN_DUMMY_13839 DFF_X1 
Xx_r3_reg_1_ n864 n6_G2B1I4 x_r3[1] NETTRAN_DUMMY_13840 NETTRAN_DUMMY_13841 NETTRAN_DUMMY_13842 DFF_X1 
Xx_r2_reg_1_ n859 n6_G2B1I4 x_r2[1] NETTRAN_DUMMY_13843 NETTRAN_DUMMY_13844 NETTRAN_DUMMY_13845 DFF_X1 
Xx_r1_reg_1_ n1840 n11_G2B1I6 x_r1[1] NETTRAN_DUMMY_13846 NETTRAN_DUMMY_13847 NETTRAN_DUMMY_13848 DFF_X1 
Xx_r3_reg_2_ n849 n10_G2B1I4 x_r3[2] NETTRAN_DUMMY_13849 NETTRAN_DUMMY_13850 NETTRAN_DUMMY_13851 DFF_X1 
Xx_r2_reg_2_ n845 n6_G2B1I2 x_r2[2] NETTRAN_DUMMY_13852 NETTRAN_DUMMY_13853 NETTRAN_DUMMY_13854 DFF_X1 
Xx_r1_reg_2_ n1820 n6_G2B1I4 x_r1[2] NETTRAN_DUMMY_13855 NETTRAN_DUMMY_13856 NETTRAN_DUMMY_13857 DFF_X1 
Xx_r3_reg_3_ n181 n6_G2B1I4 x_r3[3] NETTRAN_DUMMY_13858 NETTRAN_DUMMY_13859 NETTRAN_DUMMY_13860 DFF_X1 
Xx_r2_reg_3_ n829 n60 x_r2[3] NETTRAN_DUMMY_13861 NETTRAN_DUMMY_13862 NETTRAN_DUMMY_13863 DFF_X1 
Xx_r1_reg_3_ n180 n60_G2B1I5 x_r1[3] NETTRAN_DUMMY_13864 NETTRAN_DUMMY_13865 NETTRAN_DUMMY_13866 DFF_X1 
Xx_r3_reg_4_ n819 n10_G2B1I1 x_r3[4] NETTRAN_DUMMY_13867 NETTRAN_DUMMY_13868 NETTRAN_DUMMY_13869 DFF_X1 
Xx_r2_reg_4_ n815 n6_G2B1I2 x_r2[4] NETTRAN_DUMMY_13870 NETTRAN_DUMMY_13871 NETTRAN_DUMMY_13872 DFF_X1 
Xx_r1_reg_4_ n178 n60_G2B1I5 x_r1[4] NETTRAN_DUMMY_13873 NETTRAN_DUMMY_13874 NETTRAN_DUMMY_13875 DFF_X1 
Xx_r3_reg_5_ n804 n6_G2B1I2 x_r3[5] NETTRAN_DUMMY_13876 NETTRAN_DUMMY_13877 NETTRAN_DUMMY_13878 DFF_X1 
Xx_r2_reg_5_ n210 n6_G2B1I2 x_r2[5] NETTRAN_DUMMY_13879 NETTRAN_DUMMY_13880 NETTRAN_DUMMY_13881 DFF_X1 
Xx_r1_reg_5_ n176 n60 x_r1[5] NETTRAN_DUMMY_13882 NETTRAN_DUMMY_13883 NETTRAN_DUMMY_13884 DFF_X1 
Xx_r3_reg_6_ n789 n10_G2B1I1 x_r3[6] NETTRAN_DUMMY_13885 NETTRAN_DUMMY_13886 NETTRAN_DUMMY_13887 DFF_X1 
Xx_r2_reg_6_ n785 n10_G2B1I4 x_r2[6] NETTRAN_DUMMY_13888 NETTRAN_DUMMY_13889 NETTRAN_DUMMY_13890 DFF_X1 
Xx_r1_reg_6_ n175 n6_G2B1I4 x_r1[6] NETTRAN_DUMMY_13891 NETTRAN_DUMMY_13892 NETTRAN_DUMMY_13893 DFF_X1 
Xx_r3_reg_7_ n775 n10_G2B1I3 x_r3[7] NETTRAN_DUMMY_13894 NETTRAN_DUMMY_13895 NETTRAN_DUMMY_13896 DFF_X1 
Xsum2_rnd_reg_8_ n173 n62_G2B1I2 NETTRAN_DUMMY_13897 n35 NETTRAN_DUMMY_13898 NETTRAN_DUMMY_13899 DFF_X1 
Xsum2_rnd_reg_9_ n171 n62_G2B1I2 NETTRAN_DUMMY_13900 n34 NETTRAN_DUMMY_13901 NETTRAN_DUMMY_13902 DFF_X1 
Xsum2_rnd_reg_10_ n755 n60 NETTRAN_DUMMY_13903 n33 NETTRAN_DUMMY_13904 NETTRAN_DUMMY_13905 DFF_X1 
Xsum2_rnd_reg_11_ n170 n60_G2B1I1 NETTRAN_DUMMY_13906 n32 NETTRAN_DUMMY_13907 NETTRAN_DUMMY_13908 DFF_X1 
Xsum2_rnd_reg_12_ n169 n60_G2B1I1 NETTRAN_DUMMY_13909 n31 NETTRAN_DUMMY_13910 NETTRAN_DUMMY_13911 DFF_X1 
Xsum2_rnd_reg_13_ n168 n11_G2B1I7 NETTRAN_DUMMY_13912 n30 NETTRAN_DUMMY_13913 NETTRAN_DUMMY_13914 DFF_X1 
Xsum2_rnd_reg_14_ n167 n2 NETTRAN_DUMMY_13915 n29 NETTRAN_DUMMY_13916 NETTRAN_DUMMY_13917 DFF_X1 
Xsum2_reg_2_ N116 n7 sum2[2] NETTRAN_DUMMY_13918 NETTRAN_DUMMY_13919 NETTRAN_DUMMY_13920 DFF_X1 
Xsum2_reg_3_ N117 n7 sum2[3] NETTRAN_DUMMY_13921 NETTRAN_DUMMY_13922 NETTRAN_DUMMY_13923 DFF_X1 
Xsum2_reg_4_ N118 n9_G2B1I2 sum2[4] NETTRAN_DUMMY_13924 NETTRAN_DUMMY_13925 NETTRAN_DUMMY_13926 DFF_X1 
Xsum2_reg_5_ N119 n9_G2B1I2 sum2[5] NETTRAN_DUMMY_13927 NETTRAN_DUMMY_13928 NETTRAN_DUMMY_13929 DFF_X1 
Xsum2_reg_6_ N120 n9_G2B1I2 sum2[6] NETTRAN_DUMMY_13930 NETTRAN_DUMMY_13931 NETTRAN_DUMMY_13932 DFF_X1 
Xsum2_reg_7_ n1336 n7_G2B1I2 sum2[7] NETTRAN_DUMMY_13933 NETTRAN_DUMMY_13934 NETTRAN_DUMMY_13935 DFF_X1 
Xsum2_reg_8_ N122 n7 sum2[8] NETTRAN_DUMMY_13936 NETTRAN_DUMMY_13937 NETTRAN_DUMMY_13938 DFF_X1 
Xsum2_reg_9_ N123 n7 sum2[9] NETTRAN_DUMMY_13939 NETTRAN_DUMMY_13940 NETTRAN_DUMMY_13941 DFF_X1 
Xsum2_reg_10_ N124 n62 sum2[10] NETTRAN_DUMMY_13942 NETTRAN_DUMMY_13943 NETTRAN_DUMMY_13944 DFF_X1 
Xsum2_reg_11_ N125 n62_G2B1I2 sum2[11] NETTRAN_DUMMY_13945 NETTRAN_DUMMY_13946 NETTRAN_DUMMY_13947 DFF_X1 
Xsum2_reg_12_ N126 n63_G2B1I2 sum2[12] NETTRAN_DUMMY_13948 NETTRAN_DUMMY_13949 NETTRAN_DUMMY_13950 DFF_X1 
Xsum2_reg_13_ n1305 n60_G2B1I5 sum2[13] NETTRAN_DUMMY_13951 NETTRAN_DUMMY_13952 
+ NETTRAN_DUMMY_13953 DFF_X1 
Xsum2_reg_14_ N128 n60_G2B1I1 sum2[14] NETTRAN_DUMMY_13954 NETTRAN_DUMMY_13955 NETTRAN_DUMMY_13956 DFF_X1 
Xsum2_reg_15_ N129 n60_G2B1I1 sum2[15] NETTRAN_DUMMY_13957 NETTRAN_DUMMY_13958 NETTRAN_DUMMY_13959 DFF_X1 
Xsum2_reg_16_ N130 n11_G2B1I7 sum2[16] NETTRAN_DUMMY_13960 NETTRAN_DUMMY_13961 NETTRAN_DUMMY_13962 DFF_X1 
Xsum2_reg_17_ N131 n11_G2B1I7 NETTRAN_DUMMY_13963 n58 NETTRAN_DUMMY_13964 NETTRAN_DUMMY_13965 DFF_X1 
Xvalid_in_r_reg_8_ n732 n8_G2B1I4 valid_in_r[8] NETTRAN_DUMMY_13966 NETTRAN_DUMMY_13967 
+ NETTRAN_DUMMY_13968 DFF_X1 
Xvalid_in_r_reg_7_ n727 n8_G2B1I5 valid_in_r[7] NETTRAN_DUMMY_13969 NETTRAN_DUMMY_13970 
+ NETTRAN_DUMMY_13971 DFF_X1 
Xvalid_in_r_reg_6_ n723 n8_G2B1I8 valid_in_r[6] NETTRAN_DUMMY_13972 NETTRAN_DUMMY_13973 
+ NETTRAN_DUMMY_13974 DFF_X1 
Xvalid_in_r_reg_5_ n718 n8_G2B1I8 valid_in_r[5] NETTRAN_DUMMY_13975 NETTRAN_DUMMY_13976 
+ NETTRAN_DUMMY_13977 DFF_X1 
Xvalid_in_r_reg_4_ n714 n8_G2B1I1 valid_in_r[4] NETTRAN_DUMMY_13978 NETTRAN_DUMMY_13979 
+ NETTRAN_DUMMY_13980 DFF_X1 
Xvalid_in_r_reg_3_ n708 n8_G2B1I1 valid_in_r[3] NETTRAN_DUMMY_13981 NETTRAN_DUMMY_13982 
+ NETTRAN_DUMMY_13983 DFF_X1 
Xvalid_in_r_reg_2_ N109 n8_G2B1I7 valid_in_r[2] NETTRAN_DUMMY_13984 NETTRAN_DUMMY_13985 
+ NETTRAN_DUMMY_13986 DFF_X1 
Xvalid_in_r_reg_1_ n699 n2 valid_in_r[1] NETTRAN_DUMMY_13987 NETTRAN_DUMMY_13988 
+ NETTRAN_DUMMY_13989 DFF_X1 
Xvalid_in_r_reg_0_ n692 n2 valid_in_r[0] NETTRAN_DUMMY_13990 NETTRAN_DUMMY_13991 
+ NETTRAN_DUMMY_13992 DFF_X1 
Xsign_r_reg_8_ n691 n2 sign_r[8] n12 NETTRAN_DUMMY_13993 NETTRAN_DUMMY_13994 DFF_X1 
Xsign_r_reg_7_ n686 n2 sign_r[7] NETTRAN_DUMMY_13995 NETTRAN_DUMMY_13996 NETTRAN_DUMMY_13997 DFF_X1 
Xsign_r_reg_6_ n678 n2 sign_r[6] NETTRAN_DUMMY_13998 NETTRAN_DUMMY_13999 NETTRAN_DUMMY_14000 DFF_X1 
Xsign_r_reg_5_ n677 n2_G2B1I3 sign_r[5] NETTRAN_DUMMY_14001 NETTRAN_DUMMY_14002 
+ NETTRAN_DUMMY_14003 DFF_X1 
Xsign_r_reg_4_ n673 n2_G2B1I3 sign_r[4] NETTRAN_DUMMY_14004 NETTRAN_DUMMY_14005 
+ NETTRAN_DUMMY_14006 DFF_X1 
Xsign_r_reg_3_ n668 n2_G2B1I3 sign_r[3] NETTRAN_DUMMY_14007 NETTRAN_DUMMY_14008 
+ NETTRAN_DUMMY_14009 DFF_X1 
Xsign_r_reg_2_ n664 n2_G2B1I3 sign_r[2] NETTRAN_DUMMY_14010 NETTRAN_DUMMY_14011 
+ NETTRAN_DUMMY_14012 DFF_X1 
Xsign_r_reg_1_ n659 n2_G2B1I3 sign_r[1] NETTRAN_DUMMY_14013 NETTRAN_DUMMY_14014 
+ NETTRAN_DUMMY_14015 DFF_X1 
Xsign_r_reg_0_ data_in[0] n2_G2B1I3 sign_r[0] NETTRAN_DUMMY_14016 NETTRAN_DUMMY_14017 
+ NETTRAN_DUMMY_14018 DFF_X1 
Xc0_r5_reg_0_ n655 n8_G2B1I5 c0_r5[0] NETTRAN_DUMMY_14019 NETTRAN_DUMMY_14020 NETTRAN_DUMMY_14021 DFF_X1 
Xc0_r5_reg_1_ n651 n8_G2B1I5 c0_r5[1] NETTRAN_DUMMY_14022 NETTRAN_DUMMY_14023 NETTRAN_DUMMY_14024 DFF_X1 
Xc0_r5_reg_2_ n646 n8_G2B1I6 c0_r5[2] NETTRAN_DUMMY_14025 NETTRAN_DUMMY_14026 NETTRAN_DUMMY_14027 DFF_X1 
Xc0_r5_reg_3_ n642 n8_G2B1I6 c0_r5[3] NETTRAN_DUMMY_14028 NETTRAN_DUMMY_14029 NETTRAN_DUMMY_14030 DFF_X1 
Xc0_r5_reg_4_ n637 n7_G2B1I2 c0_r5[4] NETTRAN_DUMMY_14031 NETTRAN_DUMMY_14032 NETTRAN_DUMMY_14033 DFF_X1 
Xc0_r5_reg_5_ n633 n9_G2B1I2 c0_r5[5] NETTRAN_DUMMY_14034 NETTRAN_DUMMY_14035 NETTRAN_DUMMY_14036 DFF_X1 
Xc0_r5_reg_6_ n628 n9_G2B1I1 c0_r5[6] NETTRAN_DUMMY_14037 NETTRAN_DUMMY_14038 NETTRAN_DUMMY_14039 DFF_X1 
Xc0_r5_reg_7_ n624 n7_G2B1I1 c0_r5[7] NETTRAN_DUMMY_14040 NETTRAN_DUMMY_14041 NETTRAN_DUMMY_14042 DFF_X1 
Xc0_r5_reg_8_ n619 n7_G2B1I4 c0_r5[8] NETTRAN_DUMMY_14043 NETTRAN_DUMMY_14044 NETTRAN_DUMMY_14045 DFF_X1 
Xc0_r5_reg_9_ n615 n7_G2B1I4 c0_r5[9] NETTRAN_DUMMY_14046 NETTRAN_DUMMY_14047 NETTRAN_DUMMY_14048 DFF_X1 
Xc0_r5_reg_10_ n609 n62 c0_r5[10] NETTRAN_DUMMY_14049 NETTRAN_DUMMY_14050 NETTRAN_DUMMY_14051 DFF_X1 
Xc0_r5_reg_11_ n605 n6_G2B1I5 c0_r5[11] NETTRAN_DUMMY_14052 NETTRAN_DUMMY_14053 
+ NETTRAN_DUMMY_14054 DFF_X1 
Xc0_r5_reg_12_ n601 n6_G2B1I5 c0_r5[12] NETTRAN_DUMMY_14055 NETTRAN_DUMMY_14056 
+ NETTRAN_DUMMY_14057 DFF_X1 
Xc0_r5_reg_13_ n596 n60_G2B1I5 c0_r5[13] NETTRAN_DUMMY_14058 NETTRAN_DUMMY_14059 
+ NETTRAN_DUMMY_14060 DFF_X1 
Xc0_r5_reg_14_ n140 n2 c0_r5[14] NETTRAN_DUMMY_14061 NETTRAN_DUMMY_14062 NETTRAN_DUMMY_14063 DFF_X1 
Xc0_r5_reg_15_ n588 n11_G2B1I1 c0_r5[15] NETTRAN_DUMMY_14064 NETTRAN_DUMMY_14065 
+ NETTRAN_DUMMY_14066 DFF_X1 
Xc0_r5_reg_16_ n584 n8_G2B1I7 c0_r5[16] NETTRAN_DUMMY_14067 NETTRAN_DUMMY_14068 
+ NETTRAN_DUMMY_14069 DFF_X1 
Xc0_r5_reg_17_ n580 n11_G2B1I1 c0_r5[17] NETTRAN_DUMMY_14070 NETTRAN_DUMMY_14071 
+ NETTRAN_DUMMY_14072 DFF_X1 
Xc0_r4_reg_0_ n576 n8_G2B1I5 c0_r4[0] NETTRAN_DUMMY_14073 NETTRAN_DUMMY_14074 NETTRAN_DUMMY_14075 DFF_X1 
Xc0_r3_reg_0_ n572 n8_G2B1I5 c0_r3[0] NETTRAN_DUMMY_14076 NETTRAN_DUMMY_14077 NETTRAN_DUMMY_14078 DFF_X1 
Xc0_r2_reg_0_ n568 n8_G2B1I8 c0_r2[0] NETTRAN_DUMMY_14079 NETTRAN_DUMMY_14080 NETTRAN_DUMMY_14081 DFF_X1 
Xc0_r1_reg_0_ c0[0] n8_G2B1I8 c0_r1[0] NETTRAN_DUMMY_14082 NETTRAN_DUMMY_14083 NETTRAN_DUMMY_14084 DFF_X1 
Xc0_r4_reg_1_ n564 n8_G2B1I5 c0_r4[1] NETTRAN_DUMMY_14085 NETTRAN_DUMMY_14086 NETTRAN_DUMMY_14087 DFF_X1 
Xc0_r3_reg_1_ n560 n8_G2B1I8 c0_r3[1] NETTRAN_DUMMY_14088 NETTRAN_DUMMY_14089 NETTRAN_DUMMY_14090 DFF_X1 
Xc0_r2_reg_1_ n556 n8_G2B1I8 c0_r2[1] NETTRAN_DUMMY_14091 NETTRAN_DUMMY_14092 NETTRAN_DUMMY_14093 DFF_X1 
Xc0_r1_reg_1_ c0[1] n8_G2B1I8 c0_r1[1] NETTRAN_DUMMY_14094 NETTRAN_DUMMY_14095 NETTRAN_DUMMY_14096 DFF_X1 
Xc0_r4_reg_2_ n552 n8_G2B1I6 c0_r4[2] NETTRAN_DUMMY_14097 NETTRAN_DUMMY_14098 NETTRAN_DUMMY_14099 DFF_X1 
Xc0_r3_reg_2_ n548 n8_G2B1I6 c0_r3[2] NETTRAN_DUMMY_14100 NETTRAN_DUMMY_14101 NETTRAN_DUMMY_14102 DFF_X1 
Xc0_r2_reg_2_ n544 n8_G2B1I4 c0_r2[2] NETTRAN_DUMMY_14103 NETTRAN_DUMMY_14104 NETTRAN_DUMMY_14105 DFF_X1 
Xc0_r1_reg_2_ c0[2] n8_G2B1I4 c0_r1[2] NETTRAN_DUMMY_14106 NETTRAN_DUMMY_14107 NETTRAN_DUMMY_14108 DFF_X1 
Xc0_r4_reg_3_ n540 n8_G2B1I6 c0_r4[3] NETTRAN_DUMMY_14109 NETTRAN_DUMMY_14110 NETTRAN_DUMMY_14111 DFF_X1 
Xc0_r3_reg_3_ n536 n8_G2B1I4 c0_r3[3] NETTRAN_DUMMY_14112 NETTRAN_DUMMY_14113 NETTRAN_DUMMY_14114 DFF_X1 
Xc0_r2_reg_3_ n532 n8_G2B1I4 c0_r2[3] NETTRAN_DUMMY_14115 NETTRAN_DUMMY_14116 NETTRAN_DUMMY_14117 DFF_X1 
Xc0_r1_reg_3_ c0[3] n8_G2B1I4 c0_r1[3] NETTRAN_DUMMY_14118 NETTRAN_DUMMY_14119 NETTRAN_DUMMY_14120 DFF_X1 
Xc0_r4_reg_4_ n528 n7_G2B1I2 c0_r4[4] NETTRAN_DUMMY_14121 NETTRAN_DUMMY_14122 NETTRAN_DUMMY_14123 DFF_X1 
Xc0_r3_reg_4_ n524 n7_G2B1I2 c0_r3[4] NETTRAN_DUMMY_14124 NETTRAN_DUMMY_14125 NETTRAN_DUMMY_14126 DFF_X1 
Xc0_r2_reg_4_ n520 n7_G2B1I1 c0_r2[4] NETTRAN_DUMMY_14127 NETTRAN_DUMMY_14128 NETTRAN_DUMMY_14129 DFF_X1 
Xc0_r1_reg_4_ c0[4] n7_G2B1I1 c0_r1[4] NETTRAN_DUMMY_14130 NETTRAN_DUMMY_14131 NETTRAN_DUMMY_14132 DFF_X1 
Xc0_r4_reg_5_ n516 n9_G2B1I2 c0_r4[5] NETTRAN_DUMMY_14133 NETTRAN_DUMMY_14134 NETTRAN_DUMMY_14135 DFF_X1 
Xc0_r3_reg_5_ n512 n9_G2B1I2 c0_r3[5] NETTRAN_DUMMY_14136 NETTRAN_DUMMY_14137 NETTRAN_DUMMY_14138 DFF_X1 
Xc0_r2_reg_5_ n508 n7_G2B1I2 c0_r2[5] NETTRAN_DUMMY_14139 NETTRAN_DUMMY_14140 NETTRAN_DUMMY_14141 DFF_X1 
Xc0_r1_reg_5_ c0[5] n7_G2B1I1 c0_r1[5] NETTRAN_DUMMY_14142 NETTRAN_DUMMY_14143 NETTRAN_DUMMY_14144 DFF_X1 
Xc0_r4_reg_6_ n504 n9_G2B1I1 c0_r4[6] NETTRAN_DUMMY_14145 NETTRAN_DUMMY_14146 NETTRAN_DUMMY_14147 DFF_X1 
Xc0_r3_reg_6_ n500 n9_G2B1I1 c0_r3[6] NETTRAN_DUMMY_14148 NETTRAN_DUMMY_14149 NETTRAN_DUMMY_14150 DFF_X1 
Xc0_r2_reg_6_ n496 n9_G2B1I1 c0_r2[6] NETTRAN_DUMMY_14151 NETTRAN_DUMMY_14152 NETTRAN_DUMMY_14153 DFF_X1 
Xc0_r1_reg_6_ c0[6] n7_G2B1I2 c0_r1[6] NETTRAN_DUMMY_14154 NETTRAN_DUMMY_14155 NETTRAN_DUMMY_14156 DFF_X1 
Xc0_r4_reg_7_ n492 n8_G2B1I6 c0_r4[7] NETTRAN_DUMMY_14157 NETTRAN_DUMMY_14158 NETTRAN_DUMMY_14159 DFF_X1 
Xc0_r3_reg_7_ n488 n8_G2B1I6 c0_r3[7] NETTRAN_DUMMY_14160 NETTRAN_DUMMY_14161 NETTRAN_DUMMY_14162 DFF_X1 
Xc0_r2_reg_7_ n484 n8_G2B1I6 c0_r2[7] NETTRAN_DUMMY_14163 NETTRAN_DUMMY_14164 NETTRAN_DUMMY_14165 DFF_X1 
Xc0_r1_reg_7_ c0[7] n8_G2B1I6 c0_r1[7] NETTRAN_DUMMY_14166 NETTRAN_DUMMY_14167 NETTRAN_DUMMY_14168 DFF_X1 
Xc0_r4_reg_8_ n480 n7_G2B1I4 c0_r4[8] NETTRAN_DUMMY_14169 NETTRAN_DUMMY_14170 NETTRAN_DUMMY_14171 DFF_X1 
Xc0_r3_reg_8_ n476 n7_G2B1I4 c0_r3[8] NETTRAN_DUMMY_14172 NETTRAN_DUMMY_14173 NETTRAN_DUMMY_14174 DFF_X1 
XU71 data_in[16] rstn N78 NETTRAN_DUMMY_14175 NETTRAN_DUMMY_14176 AND2_X1 
XU70 rstn data_in[3] N91 NETTRAN_DUMMY_14177 NETTRAN_DUMMY_14178 AND2_X1 
XU69 data_in[10] rstn N84 NETTRAN_DUMMY_14179 NETTRAN_DUMMY_14180 AND2_X1 
XU68 data_in[14] rstn N80 NETTRAN_DUMMY_14181 NETTRAN_DUMMY_14182 AND2_X1 
XU67 data_in[6] rstn N88 NETTRAN_DUMMY_14183 NETTRAN_DUMMY_14184 AND2_X1 
XU66 n53 n1110 N600 NETTRAN_DUMMY_14185 NETTRAN_DUMMY_14186 NAND2_X1 
XU65 n44 n1125 n50 NETTRAN_DUMMY_14187 NETTRAN_DUMMY_14188 AND2_X1 
XU64 n1133 n7310 N611 NETTRAN_DUMMY_14189 NETTRAN_DUMMY_14190 NAND2_X1 
XU63 n1010 n910 n810 n54 NETTRAN_DUMMY_14191 NETTRAN_DUMMY_14192 NOR3_X1 
XU62 rstn n710 n6810 n54 n53 NETTRAN_DUMMY_14193 NETTRAN_DUMMY_14194 AND4_X1 
XU61 n10921 rstn n6810 n44 NETTRAN_DUMMY_14195 NETTRAN_DUMMY_14196 AND3_X1 
XU60 n7011 n1096 n44 n45 N74 NETTRAN_DUMMY_14197 NETTRAN_DUMMY_14198 NAND4_X1 
XU59 n1084 n1127 n52 NETTRAN_DUMMY_14199 NETTRAN_DUMMY_14200 AND2_X1 
XU58 n1084 n7011 n47 NETTRAN_DUMMY_14201 NETTRAN_DUMMY_14202 AND2_X1 
XU57 n44 n1127 n1096 n51 NETTRAN_DUMMY_14203 NETTRAN_DUMMY_14204 AND3_X1 
XU56 N1800 n990 NETTRAN_DUMMY_14205 NETTRAN_DUMMY_14206 INV_X1 
XU55 n55 n990 n29 n56 N196 NETTRAN_DUMMY_14207 NETTRAN_DUMMY_14208 OAI22_X1 
XU54 N1790 n1000 NETTRAN_DUMMY_14209 NETTRAN_DUMMY_14210 INV_X1 
XU53 n55 n1000 n30 n56 N195 NETTRAN_DUMMY_14211 NETTRAN_DUMMY_14212 OAI22_X1 
XU52 N1780 n1011 NETTRAN_DUMMY_14213 NETTRAN_DUMMY_14214 INV_X1 
XU51 n55 n1011 n31 n56 N194 NETTRAN_DUMMY_14215 NETTRAN_DUMMY_14216 OAI22_X1 
XU50 N1770 n1020 NETTRAN_DUMMY_14217 NETTRAN_DUMMY_14218 INV_X1 
XU49 n55 n1020 n32 n56 N193 NETTRAN_DUMMY_14219 NETTRAN_DUMMY_14220 OAI22_X1 
XU48 N1760 n1030 NETTRAN_DUMMY_14221 NETTRAN_DUMMY_14222 INV_X1 
XU47 n55 n1030 n33 n56 N192 NETTRAN_DUMMY_14223 NETTRAN_DUMMY_14224 OAI22_X1 
XU46 N1750 n1040 NETTRAN_DUMMY_14225 NETTRAN_DUMMY_14226 INV_X1 
XU45 n55 n1040 n34 n56 N191 NETTRAN_DUMMY_14227 NETTRAN_DUMMY_14228 OAI22_X1 
XU44 N1740 n1050 NETTRAN_DUMMY_14229 NETTRAN_DUMMY_14230 INV_X1 
XU43 n55 n1050 n35 n56 N190 NETTRAN_DUMMY_14231 NETTRAN_DUMMY_14232 OAI22_X1 
XU42 N1730 n1060 NETTRAN_DUMMY_14233 NETTRAN_DUMMY_14234 INV_X1 
XU41 n55 n1060 n36 n56 N189 NETTRAN_DUMMY_14235 NETTRAN_DUMMY_14236 OAI22_X1 
XU40 N1720 n1070 NETTRAN_DUMMY_14237 NETTRAN_DUMMY_14238 INV_X1 
XU39 n55 n1070 n37 n56 N188 NETTRAN_DUMMY_14239 NETTRAN_DUMMY_14240 OAI22_X1 
XU38 N1710 n1080 NETTRAN_DUMMY_14241 NETTRAN_DUMMY_14242 INV_X1 
XU37 n55 n1080 n38 n56 N187 NETTRAN_DUMMY_14243 NETTRAN_DUMMY_14244 OAI22_X1 
XU36 N1700 n1090 NETTRAN_DUMMY_14245 NETTRAN_DUMMY_14246 INV_X1 
XU35 n55 n1090 n39 n56 N186 NETTRAN_DUMMY_14247 NETTRAN_DUMMY_14248 OAI22_X1 
XU34 N1690 n1100 NETTRAN_DUMMY_14249 NETTRAN_DUMMY_14250 INV_X1 
XU33 n55 n1100 n40 n56 N185 NETTRAN_DUMMY_14251 NETTRAN_DUMMY_14252 OAI22_X1 
XU32 N1680 n1111 NETTRAN_DUMMY_14253 NETTRAN_DUMMY_14254 INV_X1 
XU31 n55 n1111 n41 n56 N184 NETTRAN_DUMMY_14255 NETTRAN_DUMMY_14256 OAI22_X1 
XU30 N1670 n1120 NETTRAN_DUMMY_14257 NETTRAN_DUMMY_14258 INV_X1 
XU29 n55 n1120 n42 n56 N183 NETTRAN_DUMMY_14259 NETTRAN_DUMMY_14260 OAI22_X1 
XU28 n55 n43 n43 n56 N182 NETTRAN_DUMMY_14261 NETTRAN_DUMMY_14262 OAI22_X1 
XU25 rstn n12 n56 NETTRAN_DUMMY_14263 NETTRAN_DUMMY_14264 NAND2_X1 
XU24 sign_r[8] rstn n55 NETTRAN_DUMMY_14265 NETTRAN_DUMMY_14266 NAND2_X1 
XU23 num_lzd[5] rstn N11000 NETTRAN_DUMMY_14267 NETTRAN_DUMMY_14268 AND2_X1 
XU22 num_lzd[4] rstn N10 NETTRAN_DUMMY_14269 NETTRAN_DUMMY_14270 AND2_X1 
XU21 num_lzd[2] rstn N8 NETTRAN_DUMMY_14271 NETTRAN_DUMMY_14272 AND2_X1 
XU20 num_lzd[3] rstn N900 NETTRAN_DUMMY_14273 NETTRAN_DUMMY_14274 AND2_X1 
XU19 num_lzd[1] rstn N700 NETTRAN_DUMMY_14275 NETTRAN_DUMMY_14276 AND2_X1 
XU18 num_lzd[0] rstn N610 NETTRAN_DUMMY_14277 NETTRAN_DUMMY_14278 AND2_X1 
XU17 n52 n1107 N65 NETTRAN_DUMMY_14279 NETTRAN_DUMMY_14280 NAND2_X1 
XU16 n52 n1115 N64 NETTRAN_DUMMY_14281 NETTRAN_DUMMY_14282 NAND2_X1 
XU15 n52 n1119 N63 NETTRAN_DUMMY_14283 NETTRAN_DUMMY_14284 NAND2_X1 
XU14 n51 n1107 N69 NETTRAN_DUMMY_14285 NETTRAN_DUMMY_14286 NAND2_X1 
XU13 n51 n1115 N68 NETTRAN_DUMMY_14287 NETTRAN_DUMMY_14288 NAND2_X1 
XU12 n51 n1119 N67 NETTRAN_DUMMY_14289 NETTRAN_DUMMY_14290 NAND2_X1 
XU11 n47 n45 N7010 NETTRAN_DUMMY_14291 NETTRAN_DUMMY_14292 NAND2_X1 
XU10 n51 n45 N66 NETTRAN_DUMMY_14293 NETTRAN_DUMMY_14294 NAND2_X1 
XU9 n52 n45 N620 NETTRAN_DUMMY_14295 NETTRAN_DUMMY_14296 NAND2_X1 
XU8 n1107 n47 N73 NETTRAN_DUMMY_14297 NETTRAN_DUMMY_14298 NAND2_X1 
XU6 n1115 n47 N72 NETTRAN_DUMMY_14299 NETTRAN_DUMMY_14300 NAND2_X1 
XU5 n1119 n47 N71 NETTRAN_DUMMY_14301 NETTRAN_DUMMY_14302 NAND2_X1 
XU4 N1810 n980 NETTRAN_DUMMY_14303 NETTRAN_DUMMY_14304 INV_X1 
XU3 n980 n55 N197 NETTRAN_DUMMY_14305 NETTRAN_DUMMY_14306 NOR2_X1 
Xdata_out_reg_0_ n166 n9_G2B1I1 data_out[0] NETTRAN_DUMMY_14307 NETTRAN_DUMMY_14308 
+ NETTRAN_DUMMY_14309 DFF_X1 
Xdata_out_reg_1_ n462 n9_G2B1I2 data_out[1] NETTRAN_DUMMY_14310 NETTRAN_DUMMY_14311 
+ NETTRAN_DUMMY_14312 DFF_X1 
Xdata_out_reg_2_ n456 n7_G2B1I1 data_out[2] NETTRAN_DUMMY_14313 NETTRAN_DUMMY_14314 
+ NETTRAN_DUMMY_14315 DFF_X1 
Xdata_out_reg_3_ n139 clk_G1B1I5 data_out[3] NETTRAN_DUMMY_14316 NETTRAN_DUMMY_14317 
+ NETTRAN_DUMMY_14318 DFF_X1 
Xdata_out_reg_4_ n1304 n8_G2B1I4 data_out[4] NETTRAN_DUMMY_14319 NETTRAN_DUMMY_14320 
+ NETTRAN_DUMMY_14321 DFF_X1 
Xdata_out_reg_5_ n165 n61_G2B1I1 data_out[5] NETTRAN_DUMMY_14322 NETTRAN_DUMMY_14323 
+ NETTRAN_DUMMY_14324 DFF_X1 
Xdata_out_reg_6_ n164 n61_G2B1I1 data_out[6] NETTRAN_DUMMY_14325 NETTRAN_DUMMY_14326 
+ NETTRAN_DUMMY_14327 DFF_X1 
Xdata_out_reg_7_ n138 n61_G2B1I1 data_out[7] NETTRAN_DUMMY_14328 NETTRAN_DUMMY_14329 
+ NETTRAN_DUMMY_14330 DFF_X1 
Xdata_out_reg_8_ n1333 n9_G2B1I1 data_out[8] NETTRAN_DUMMY_14331 NETTRAN_DUMMY_14332 
+ NETTRAN_DUMMY_14333 DFF_X1 
Xdata_out_reg_9_ n420 n9_G2B1I1 data_out[9] NETTRAN_DUMMY_14334 NETTRAN_DUMMY_14335 
+ NETTRAN_DUMMY_14336 DFF_X1 
Xdata_out_reg_10_ n137 n60 data_out[10] NETTRAN_DUMMY_14337 NETTRAN_DUMMY_14338 
+ NETTRAN_DUMMY_14339 DFF_X1 
Xdata_out_reg_11_ n408 n60 data_out[11] NETTRAN_DUMMY_14340 NETTRAN_DUMMY_14341 
+ NETTRAN_DUMMY_14342 DFF_X1 
Xdata_out_reg_12_ n162 n60_G2B1I1 data_out[12] NETTRAN_DUMMY_14343 NETTRAN_DUMMY_14344 
+ NETTRAN_DUMMY_14345 DFF_X1 
Xdata_out_reg_13_ n400 n2 data_out[13] NETTRAN_DUMMY_14346 NETTRAN_DUMMY_14347 NETTRAN_DUMMY_14348 DFF_X1 
Xdata_out_reg_14_ n136 n2_G2B1I3 data_out[14] NETTRAN_DUMMY_14349 NETTRAN_DUMMY_14350 
+ NETTRAN_DUMMY_14351 DFF_X1 
Xdata_out_reg_15_ n160 n2_G2B1I3 data_out[15] NETTRAN_DUMMY_14352 NETTRAN_DUMMY_14353 
+ NETTRAN_DUMMY_14354 DFF_X1 
Xvalid_out_reg n386 n8_G2B1I4 valid_out NETTRAN_DUMMY_14355 NETTRAN_DUMMY_14356 
+ NETTRAN_DUMMY_14357 DFF_X1 
Xsum2_rnd_reg_0_ n158 n7 NETTRAN_DUMMY_14358 n43 NETTRAN_DUMMY_14359 NETTRAN_DUMMY_14360 DFF_X1 
Xsum2_rnd_reg_1_ n157 n9_G2B1I2 NETTRAN_DUMMY_14361 n42 NETTRAN_DUMMY_14362 NETTRAN_DUMMY_14363 DFF_X1 
Xsum2_rnd_reg_2_ n156 n9_G2B1I2 NETTRAN_DUMMY_14364 n41 NETTRAN_DUMMY_14365 NETTRAN_DUMMY_14366 DFF_X1 
Xsum2_rnd_reg_3_ n155 n9_G2B1I2 NETTRAN_DUMMY_14367 n40 NETTRAN_DUMMY_14368 NETTRAN_DUMMY_14369 DFF_X1 
Xsum2_rnd_reg_4_ n154 n7_G2B1I2 NETTRAN_DUMMY_14370 n39 NETTRAN_DUMMY_14371 NETTRAN_DUMMY_14372 DFF_X1 
Xsum2_rnd_reg_5_ n153 n7 NETTRAN_DUMMY_14373 n38 NETTRAN_DUMMY_14374 NETTRAN_DUMMY_14375 DFF_X1 
Xsum2_rnd_reg_6_ n152 n7 NETTRAN_DUMMY_14376 n37 NETTRAN_DUMMY_14377 NETTRAN_DUMMY_14378 DFF_X1 
Xsum2_rnd_reg_7_ n151 n62 NETTRAN_DUMMY_14379 n36 NETTRAN_DUMMY_14380 NETTRAN_DUMMY_14381 DFF_X1 
XU141 sum2[8] n5 n940 NETTRAN_DUMMY_14382 NETTRAN_DUMMY_14383 XOR2_X1 
XU140 sum2[7] n17 n930 NETTRAN_DUMMY_14384 NETTRAN_DUMMY_14385 XOR2_X1 
XU139 sum2[6] n16 n920 NETTRAN_DUMMY_14386 NETTRAN_DUMMY_14387 XOR2_X1 
XU138 sum2[5] n4 n911 NETTRAN_DUMMY_14388 NETTRAN_DUMMY_14389 XOR2_X1 
XU137 sum2[4] n3 n9000 NETTRAN_DUMMY_14390 NETTRAN_DUMMY_14391 XOR2_X1 
XU136 sum2[2] sum2[3] n890 NETTRAN_DUMMY_14392 NETTRAN_DUMMY_14393 XOR2_X1 
XU135 n870 n880 N92 NETTRAN_DUMMY_14394 NETTRAN_DUMMY_14395 NOR2_X1 
XU134 n850 n860 N93 NETTRAN_DUMMY_14396 NETTRAN_DUMMY_14397 NOR2_X1 
XU133 n830 n840 N94 NETTRAN_DUMMY_14398 NETTRAN_DUMMY_14399 NOR2_X1 
XU132 n811 n820 N95 NETTRAN_DUMMY_14400 NETTRAN_DUMMY_14401 NOR2_X1 
XU131 n790 n800 N96 NETTRAN_DUMMY_14402 NETTRAN_DUMMY_14403 NOR2_X1 
XU130 n770 n780 N97 NETTRAN_DUMMY_14404 NETTRAN_DUMMY_14405 NOR2_X1 
XU129 n750 n760 N98 NETTRAN_DUMMY_14406 NETTRAN_DUMMY_14407 NOR2_X1 
XU128 n730 n740 N99 NETTRAN_DUMMY_14408 NETTRAN_DUMMY_14409 NOR2_X1 
XU127 n711 n720 N100 NETTRAN_DUMMY_14410 NETTRAN_DUMMY_14411 NOR2_X1 
XU126 n690 n7000 N101 NETTRAN_DUMMY_14412 NETTRAN_DUMMY_14413 NOR2_X1 
XU125 n670 n680 N102 NETTRAN_DUMMY_14414 NETTRAN_DUMMY_14415 NOR2_X1 
XU124 n650 n660 N103 NETTRAN_DUMMY_14416 NETTRAN_DUMMY_14417 NOR2_X1 
XU123 n630 n640 N104 NETTRAN_DUMMY_14418 NETTRAN_DUMMY_14419 NOR2_X1 
XU122 n6110 n6200 N105 NETTRAN_DUMMY_14420 NETTRAN_DUMMY_14421 NOR2_X1 
XU121 n59 n6000 N106 NETTRAN_DUMMY_14422 NETTRAN_DUMMY_14423 NOR2_X1 
XU120 n1091 n1095 n46 NETTRAN_DUMMY_14424 NETTRAN_DUMMY_14425 NOR2_X1 
XU119 n1091 n7310 n48 NETTRAN_DUMMY_14426 NETTRAN_DUMMY_14427 NOR2_X1 
XU118 n1095 n7210 n49 NETTRAN_DUMMY_14428 NETTRAN_DUMMY_14429 NOR2_X1 
XU117 n1086 n7310 n45 NETTRAN_DUMMY_14430 NETTRAN_DUMMY_14431 NOR2_X1 
XU116 sum2[16] n15 n950 NETTRAN_DUMMY_14432 NETTRAN_DUMMY_14433 NAND2_X1 
XU115 n58 n950 n57 NETTRAN_DUMMY_14434 NETTRAN_DUMMY_14435 XOR2_X1 
XU114 sum2[16] n15 n28 NETTRAN_DUMMY_14436 NETTRAN_DUMMY_14437 XOR2_X1 
XU113 sum2[15] n21 n27 NETTRAN_DUMMY_14438 NETTRAN_DUMMY_14439 XOR2_X1 
XU112 sum2[14] n20 n26 NETTRAN_DUMMY_14440 NETTRAN_DUMMY_14441 XOR2_X1 
XU111 sum2[13] n14 n25 NETTRAN_DUMMY_14442 NETTRAN_DUMMY_14443 XOR2_X1 
XU110 sum2[12] n19 n24 NETTRAN_DUMMY_14444 NETTRAN_DUMMY_14445 XOR2_X1 
XU109 sum2[11] n18 n23 NETTRAN_DUMMY_14446 NETTRAN_DUMMY_14447 XOR2_X1 
XU108 sum2[10] n13 n22 NETTRAN_DUMMY_14448 NETTRAN_DUMMY_14449 XOR2_X1 
XU107 sum2[14] n20 n21 NETTRAN_DUMMY_14450 NETTRAN_DUMMY_14451 AND2_X1 
XU106 sum2[13] n14 n20 NETTRAN_DUMMY_14452 NETTRAN_DUMMY_14453 AND2_X1 
XU105 sum2[11] n18 n19 NETTRAN_DUMMY_14454 NETTRAN_DUMMY_14455 AND2_X1 
XU104 sum2[10] n13 n18 NETTRAN_DUMMY_14456 NETTRAN_DUMMY_14457 AND2_X1 
XU103 sum2[6] n16 n17 NETTRAN_DUMMY_14458 NETTRAN_DUMMY_14459 AND2_X1 
XU102 sum2[5] n4 n16 NETTRAN_DUMMY_14460 NETTRAN_DUMMY_14461 AND2_X1 
XU101 sum2[15] n21 n15 NETTRAN_DUMMY_14462 NETTRAN_DUMMY_14463 AND2_X1 
XU100 sum2[12] n19 n14 NETTRAN_DUMMY_14464 NETTRAN_DUMMY_14465 AND2_X1 
XU99 sum2[9] n6100 n13 NETTRAN_DUMMY_14466 NETTRAN_DUMMY_14467 AND2_X1 
XU98 sum2[8] n5 n6100 NETTRAN_DUMMY_14468 NETTRAN_DUMMY_14469 AND2_X1 
XU97 sum2[7] n17 n5 NETTRAN_DUMMY_14470 NETTRAN_DUMMY_14471 AND2_X1 
XU96 sum2[4] n3 n4 NETTRAN_DUMMY_14472 NETTRAN_DUMMY_14473 AND2_X1 
XU95 sum2[2] sum2[3] n3 NETTRAN_DUMMY_14474 NETTRAN_DUMMY_14475 AND2_X1 
XU94 sum2[9] n6100 n1 NETTRAN_DUMMY_14476 NETTRAN_DUMMY_14477 XOR2_X1 
XU93 data_in[1] IN1 N76 NETTRAN_DUMMY_14478 NETTRAN_DUMMY_14479 AND2_X1 
XU92 data_in[2] IN0 N75 NETTRAN_DUMMY_14480 NETTRAN_DUMMY_14481 AND2_X1 
XU91 data_in[17] rstn N77 NETTRAN_DUMMY_14482 NETTRAN_DUMMY_14483 AND2_X1 
XU90 valid_in IN2 N107 NETTRAN_DUMMY_14484 NETTRAN_DUMMY_14485 AND2_X1 
XU89 valid_in_r[0] IN2 N108 NETTRAN_DUMMY_14486 NETTRAN_DUMMY_14487 AND2_X1 
XU88 n704 IN1 N109 NETTRAN_DUMMY_14488 NETTRAN_DUMMY_14489 AND2_X1 
XU87 valid_in_r[2] IN1 N11010 NETTRAN_DUMMY_14490 NETTRAN_DUMMY_14491 AND2_X1 
XU86 valid_in_r[3] IN1 N111 NETTRAN_DUMMY_14492 NETTRAN_DUMMY_14493 AND2_X1 
XU85 valid_in_r[4] IN1 N112 NETTRAN_DUMMY_14494 NETTRAN_DUMMY_14495 AND2_X1 
XU84 valid_in_r[5] IN1 N113 NETTRAN_DUMMY_14496 NETTRAN_DUMMY_14497 AND2_X1 
XU83 valid_in_r[6] IN1 N114 NETTRAN_DUMMY_14498 NETTRAN_DUMMY_14499 AND2_X1 
XU82 valid_in_r[7] IN1 N115 NETTRAN_DUMMY_14500 NETTRAN_DUMMY_14501 AND2_X1 
XU81 valid_in_r[8] IN1 N147 NETTRAN_DUMMY_14502 NETTRAN_DUMMY_14503 AND2_X1 
XU80 data_in[4] rstn N9010 NETTRAN_DUMMY_14504 NETTRAN_DUMMY_14505 AND2_X1 
XU79 data_in[5] rstn N89 NETTRAN_DUMMY_14506 NETTRAN_DUMMY_14507 AND2_X1 
XU78 data_in[7] rstn N87 NETTRAN_DUMMY_14508 NETTRAN_DUMMY_14509 AND2_X1 
XU77 data_in[8] rstn N86 NETTRAN_DUMMY_14510 NETTRAN_DUMMY_14511 AND2_X1 
XU76 data_in[9] rstn N85 NETTRAN_DUMMY_14512 NETTRAN_DUMMY_14513 AND2_X1 
XU75 data_in[11] rstn N83 NETTRAN_DUMMY_14514 NETTRAN_DUMMY_14515 AND2_X1 
XU74 data_in[12] rstn N82 NETTRAN_DUMMY_14516 NETTRAN_DUMMY_14517 AND2_X1 
XU73 data_in[13] rstn N81 NETTRAN_DUMMY_14518 NETTRAN_DUMMY_14519 AND2_X1 
XU72 data_in[15] rstn N79 NETTRAN_DUMMY_14520 NETTRAN_DUMMY_14521 AND2_X1 
XU145 clk_G1B1I7 n6111 NETTRAN_DUMMY_14522 NETTRAN_DUMMY_14523 BUF_X32 
XU142 clk_G1B1I7 n10920 NETTRAN_DUMMY_14524 NETTRAN_DUMMY_14525 BUF_X32 
XCLKBUF_X1_G2B1I1 n11 n11_G2B1I1 NETTRAN_DUMMY_14526 NETTRAN_DUMMY_14527 CLKBUF_X1 
XCLKBUF_X1_G2B1I2 n11 n11_G2B1I2 NETTRAN_DUMMY_14528 NETTRAN_DUMMY_14529 CLKBUF_X1 
XCLKBUF_X1_G2B1I3 n11 n11_G2B1I3 NETTRAN_DUMMY_14530 NETTRAN_DUMMY_14531 CLKBUF_X1 
XCLKBUF_X1_G2B1I4 n11 n11_G2B1I4 NETTRAN_DUMMY_14532 NETTRAN_DUMMY_14533 CLKBUF_X1 
XCLKBUF_X1_G2B1I5 n11 n11_G2B1I5 NETTRAN_DUMMY_14534 NETTRAN_DUMMY_14535 CLKBUF_X1 
XCLKBUF_X1_G2B1I6 n11 n11_G2B1I6 NETTRAN_DUMMY_14536 NETTRAN_DUMMY_14537 CLKBUF_X1 
XCLKBUF_X1_G2B1I7 n11 n11_G2B1I7 NETTRAN_DUMMY_14538 NETTRAN_DUMMY_14539 CLKBUF_X1 
XCLKBUF_X1_G2B1I31 n2 n2_G2B1I3 NETTRAN_DUMMY_14540 NETTRAN_DUMMY_14541 CLKBUF_X1 
XCLKBUF_X1_G2B1I13 n10920 n10_G2B1I1 NETTRAN_DUMMY_14542 NETTRAN_DUMMY_14543 CLKBUF_X1 
XCLKBUF_X1_G2B1I23 n10920 n10_G2B1I2 NETTRAN_DUMMY_14544 NETTRAN_DUMMY_14545 CLKBUF_X1 
XCLKBUF_X1_G2B1I33 n10920 n10_G2B1I3 NETTRAN_DUMMY_14546 NETTRAN_DUMMY_14547 CLKBUF_X1 
XCLKBUF_X1_G2B1I42 n10920 n10_G2B1I4 NETTRAN_DUMMY_14548 NETTRAN_DUMMY_14549 CLKBUF_X1 
XCLKBUF_X1_G2B1I25 n6310 n63_G2B1I2 NETTRAN_DUMMY_14550 NETTRAN_DUMMY_14551 CLKBUF_X1 
XCLKBUF_X1_G2B1I15 clk_G1B1I5 n8_G2B1I1 NETTRAN_DUMMY_14552 NETTRAN_DUMMY_14553 CLKBUF_X1 
XCLKBUF_X1_G2B1I26 clk_G1B1I5 n8_G2B1I2 NETTRAN_DUMMY_14554 NETTRAN_DUMMY_14555 CLKBUF_X1 
XCLKBUF_X1_G2B1I44 clk_G1B1I5 n8_G2B1I4 NETTRAN_DUMMY_14556 NETTRAN_DUMMY_14557 CLKBUF_X1 
XCLKBUF_X1_G2B1I53 clk_G1B1I5 n8_G2B1I5 NETTRAN_DUMMY_14558 NETTRAN_DUMMY_14559 CLKBUF_X1 
XCLKBUF_X1_G2B1I61 clk_G1B1I5 n8_G2B1I6 NETTRAN_DUMMY_14560 NETTRAN_DUMMY_14561 CLKBUF_X1 
XCLKBUF_X1_G2B1I71 clk_G1B1I5 n8_G2B1I7 NETTRAN_DUMMY_14562 NETTRAN_DUMMY_14563 CLKBUF_X1 
XCLKBUF_X1_G2B1I81 clk_G1B1I5 n8_G2B1I8 NETTRAN_DUMMY_14564 NETTRAN_DUMMY_14565 CLKBUF_X1 
XCLKBUF_X1_G2B1I16 n7 n7_G2B1I1 NETTRAN_DUMMY_14566 NETTRAN_DUMMY_14567 CLKBUF_X1 
XCLKBUF_X1_G2B1I27 n7 n7_G2B1I2 NETTRAN_DUMMY_14568 NETTRAN_DUMMY_14569 CLKBUF_X1 
XCLKBUF_X1_G2B1I45 n7 n7_G2B1I4 NETTRAN_DUMMY_14570 NETTRAN_DUMMY_14571 CLKBUF_X1 
XCLKBUF_X1_G2B1I29 n62 n62_G2B1I2 NETTRAN_DUMMY_14572 NETTRAN_DUMMY_14573 CLKBUF_X1 
XCLKBUF_X1_G2B1I19 n6111 n61_G2B1I1 NETTRAN_DUMMY_14574 NETTRAN_DUMMY_14575 CLKBUF_X1 
XCLKBUF_X3_G1B1I7 clk clk_G1B1I7 NETTRAN_DUMMY_14576 NETTRAN_DUMMY_14577 CLKBUF_X3 
XCLKBUF_X3_G1B1I8 clk clk_G1B1I8 NETTRAN_DUMMY_14578 NETTRAN_DUMMY_14579 CLKBUF_X1 
XCLKBUF_X2_G1B1I5 clk clk_G1B1I5 NETTRAN_DUMMY_14580 NETTRAN_DUMMY_14581 CLKBUF_X1 
XCLKBUF_X3_G1B1I4 clk clk_G1B1I4 NETTRAN_DUMMY_14582 NETTRAN_DUMMY_14583 CLKBUF_X1 
XU146 clk_G1B1I4 n62 NETTRAN_DUMMY_14584 NETTRAN_DUMMY_14585 CLKBUF_X1 
XU27 clk_G1B1I4 n9 NETTRAN_DUMMY_14586 NETTRAN_DUMMY_14587 CLKBUF_X1 
XCLKBUF_X2_G1B1I1 clk clk_G1B1I1 NETTRAN_DUMMY_14588 NETTRAN_DUMMY_14589 CLKBUF_X1 
XU1 clk_cts_3 n2 NETTRAN_DUMMY_14590 NETTRAN_DUMMY_14591 CLKBUF_X1 
XU143 clk_cts_3 n11 NETTRAN_DUMMY_14592 NETTRAN_DUMMY_14593 CLKBUF_X1 
XCLKBUF_X1_G2B1I8 n6310 n63_G2B1I8 NETTRAN_DUMMY_14594 NETTRAN_DUMMY_14595 CLKBUF_X1 
XU7 clk_G1B1I4 n7 NETTRAN_DUMMY_14596 NETTRAN_DUMMY_14597 CLKBUF_X1 
XCLKBUF_X1_G2B1I17 n9 n9_G2B1I1 NETTRAN_DUMMY_14598 NETTRAN_DUMMY_14599 CLKBUF_X1 
XCLKBUF_X1_G2B1I28 n9 n9_G2B1I2 NETTRAN_DUMMY_14600 NETTRAN_DUMMY_14601 CLKBUF_X1 
XCLKBUF_X1_G2B1I22 n6 n6_G2B1I2 NETTRAN_DUMMY_14602 NETTRAN_DUMMY_14603 CLKBUF_X1 
XCLKBUF_X1_G2B1I32 n6 n6_G2B1I3 NETTRAN_DUMMY_14604 NETTRAN_DUMMY_14605 CLKBUF_X1 
XCLKBUF_X1_G2B1I41 n6 n6_G2B1I4 NETTRAN_DUMMY_14606 NETTRAN_DUMMY_14607 CLKBUF_X1 
XCLKBUF_X1_G2B1I51 n6 n6_G2B1I5 NETTRAN_DUMMY_14608 NETTRAN_DUMMY_14609 CLKBUF_X1 
XU2 clk_G1B1I8 n6 NETTRAN_DUMMY_14610 NETTRAN_DUMMY_14611 CLKBUF_X1 
XCLKBUF_X1_G2B1I14 n60 n60_G2B1I1 NETTRAN_DUMMY_14612 NETTRAN_DUMMY_14613 CLKBUF_X1 
XCLKBUF_X1_G2B1I52 n60 n60_G2B1I5 NETTRAN_DUMMY_14614 NETTRAN_DUMMY_14615 CLKBUF_X1 
XU144 clk_G1B1I8 n60 NETTRAN_DUMMY_14616 NETTRAN_DUMMY_14617 CLKBUF_X1 
XU147 clk_G1B1I1 n6310 NETTRAN_DUMMY_14618 NETTRAN_DUMMY_14619 CLKBUF_X3 
XU26 num_lzd_r[0] n132 NETTRAN_DUMMY_14620 NETTRAN_DUMMY_14621 CLKBUF_X2 
XU149 n204 n133 NETTRAN_DUMMY_14622 NETTRAN_DUMMY_14623 BUF_X1 
XU151 n1101 n134 NETTRAN_DUMMY_14624 NETTRAN_DUMMY_14625 BUF_X1 
XU154 n208 n135 NETTRAN_DUMMY_14626 NETTRAN_DUMMY_14627 BUF_X1 
XU155 n161 n136 NETTRAN_DUMMY_14628 NETTRAN_DUMMY_14629 BUF_X1 
XU156 n415 n137 NETTRAN_DUMMY_14630 NETTRAN_DUMMY_14631 BUF_X1 
XU157 n163 n138 NETTRAN_DUMMY_14632 NETTRAN_DUMMY_14633 BUF_X1 
XU158 n452 n139 NETTRAN_DUMMY_14634 NETTRAN_DUMMY_14635 BUF_X1 
XU159 n589 n140 NETTRAN_DUMMY_14636 NETTRAN_DUMMY_14637 BUF_X1 
XU160 n866 n141 NETTRAN_DUMMY_14638 NETTRAN_DUMMY_14639 BUF_X1 
XU161 n1088 n142 NETTRAN_DUMMY_14640 NETTRAN_DUMMY_14641 BUF_X1 
XU162 num_lzd_r[2] n143 NETTRAN_DUMMY_14642 NETTRAN_DUMMY_14643 BUF_X1 
XU163 n1123 n1127 NETTRAN_DUMMY_14644 NETTRAN_DUMMY_14645 INV_X16 
XU164 n1116 n1117 NETTRAN_DUMMY_14646 NETTRAN_DUMMY_14647 INV_X8 
XU165 n1108 n1109 NETTRAN_DUMMY_14648 NETTRAN_DUMMY_14649 INV_X1 
XU166 n1102 n1103 NETTRAN_DUMMY_14650 NETTRAN_DUMMY_14651 INV_X1 
XU167 n1890 n1900 NETTRAN_DUMMY_14652 NETTRAN_DUMMY_14653 INV_X1 
XU168 n144 n145 NETTRAN_DUMMY_14654 NETTRAN_DUMMY_14655 INV_X4 
XU169 n146 n1470 NETTRAN_DUMMY_14656 NETTRAN_DUMMY_14657 INV_X4 
XU170 n149 n150 NETTRAN_DUMMY_14658 NETTRAN_DUMMY_14659 INV_X1 
XU171 n238 n144 NETTRAN_DUMMY_14660 NETTRAN_DUMMY_14661 INV_X1 
XU172 n254 n146 NETTRAN_DUMMY_14662 NETTRAN_DUMMY_14663 INV_X1 
XU173 n274 n148 NETTRAN_DUMMY_14664 NETTRAN_DUMMY_14665 BUF_X1 
XU174 n273 n149 NETTRAN_DUMMY_14666 NETTRAN_DUMMY_14667 INV_X1 
XU175 n347 n151 NETTRAN_DUMMY_14668 NETTRAN_DUMMY_14669 BUF_X1 
XU176 n350 n152 NETTRAN_DUMMY_14670 NETTRAN_DUMMY_14671 BUF_X1 
XU177 n357 n153 NETTRAN_DUMMY_14672 NETTRAN_DUMMY_14673 BUF_X1 
XU178 n362 n154 NETTRAN_DUMMY_14674 NETTRAN_DUMMY_14675 BUF_X1 
XU179 n367 n155 NETTRAN_DUMMY_14676 NETTRAN_DUMMY_14677 BUF_X1 
XU180 n372 n156 NETTRAN_DUMMY_14678 NETTRAN_DUMMY_14679 BUF_X1 
XU181 n377 n157 NETTRAN_DUMMY_14680 NETTRAN_DUMMY_14681 BUF_X1 
XU182 n382 n158 NETTRAN_DUMMY_14682 NETTRAN_DUMMY_14683 BUF_X1 
XU183 n389 n159 NETTRAN_DUMMY_14684 NETTRAN_DUMMY_14685 INV_X1 
XU184 n159 n160 NETTRAN_DUMMY_14686 NETTRAN_DUMMY_14687 INV_X8 
XU185 n395 n161 NETTRAN_DUMMY_14688 NETTRAN_DUMMY_14689 CLKBUF_X1 
XU186 n407 n162 NETTRAN_DUMMY_14690 NETTRAN_DUMMY_14691 BUF_X1 
XU187 n431 n163 NETTRAN_DUMMY_14692 NETTRAN_DUMMY_14693 CLKBUF_X1 
XU188 n437 n164 NETTRAN_DUMMY_14694 NETTRAN_DUMMY_14695 BUF_X1 
XU189 n443 n165 NETTRAN_DUMMY_14696 NETTRAN_DUMMY_14697 BUF_X1 
XU190 n470 n166 NETTRAN_DUMMY_14698 NETTRAN_DUMMY_14699 BUF_X1 
XU191 n737 n167 NETTRAN_DUMMY_14700 NETTRAN_DUMMY_14701 BUF_X1 
XU192 n743 n168 NETTRAN_DUMMY_14702 NETTRAN_DUMMY_14703 BUF_X1 
XU193 n748 n169 NETTRAN_DUMMY_14704 NETTRAN_DUMMY_14705 BUF_X1 
XU194 n754 n170 NETTRAN_DUMMY_14706 NETTRAN_DUMMY_14707 BUF_X1 
XU195 n765 n171 NETTRAN_DUMMY_14708 NETTRAN_DUMMY_14709 CLKBUF_X1 
XU196 n771 n172 NETTRAN_DUMMY_14710 NETTRAN_DUMMY_14711 INV_X1 
XU197 n172 n173 NETTRAN_DUMMY_14712 NETTRAN_DUMMY_14713 INV_X8 
XU198 n778 n174 NETTRAN_DUMMY_14714 NETTRAN_DUMMY_14715 INV_X1 
XU199 n174 n175 NETTRAN_DUMMY_14716 NETTRAN_DUMMY_14717 INV_X16 
XU200 n795 n176 NETTRAN_DUMMY_14718 NETTRAN_DUMMY_14719 BUF_X1 
XU201 n809 n177 NETTRAN_DUMMY_14720 NETTRAN_DUMMY_14721 INV_X1 
XU202 n177 n178 NETTRAN_DUMMY_14722 NETTRAN_DUMMY_14723 INV_X16 
XU203 n825 n179 NETTRAN_DUMMY_14724 NETTRAN_DUMMY_14725 INV_X1 
XU204 n179 n180 NETTRAN_DUMMY_14726 NETTRAN_DUMMY_14727 INV_X16 
XU205 n834 n181 NETTRAN_DUMMY_14728 NETTRAN_DUMMY_14729 BUF_X1 
XU206 n838 n1820 NETTRAN_DUMMY_14730 NETTRAN_DUMMY_14731 BUF_X1 
XU207 n855 n1830 NETTRAN_DUMMY_14732 NETTRAN_DUMMY_14733 INV_X1 
XU208 n1830 n1840 NETTRAN_DUMMY_14734 NETTRAN_DUMMY_14735 INV_X16 
XU209 n921 n1850 NETTRAN_DUMMY_14736 NETTRAN_DUMMY_14737 BUF_X1 
XU210 n929 n1860 NETTRAN_DUMMY_14738 NETTRAN_DUMMY_14739 BUF_X1 
XU211 n1017 n1870 NETTRAN_DUMMY_14740 NETTRAN_DUMMY_14741 CLKBUF_X1 
XU212 n1057 n1880 NETTRAN_DUMMY_14742 NETTRAN_DUMMY_14743 BUF_X1 
XU213 n1056 n1890 NETTRAN_DUMMY_14744 NETTRAN_DUMMY_14745 INV_X1 
XU214 N610 n1910 NETTRAN_DUMMY_14746 NETTRAN_DUMMY_14747 INV_X1 
XU215 n1910 n1920 NETTRAN_DUMMY_14748 NETTRAN_DUMMY_14749 INV_X16 
XU216 n1158 n1930 NETTRAN_DUMMY_14750 NETTRAN_DUMMY_14751 CLKBUF_X1 
XU217 n1202 n1940 NETTRAN_DUMMY_14752 NETTRAN_DUMMY_14753 BUF_X1 
XU218 n1216 n1950 NETTRAN_DUMMY_14754 NETTRAN_DUMMY_14755 BUF_X1 
XU219 n1229 n1960 NETTRAN_DUMMY_14756 NETTRAN_DUMMY_14757 INV_X1 
XU220 n1960 n1970 NETTRAN_DUMMY_14758 NETTRAN_DUMMY_14759 INV_X16 
XU221 n1245 n198 NETTRAN_DUMMY_14760 NETTRAN_DUMMY_14761 BUF_X1 
XU222 n1258 n199 NETTRAN_DUMMY_14762 NETTRAN_DUMMY_14763 INV_X1 
XU223 n199 n200 NETTRAN_DUMMY_14764 NETTRAN_DUMMY_14765 INV_X16 
XU224 n1299 n201 NETTRAN_DUMMY_14766 NETTRAN_DUMMY_14767 BUF_X1 
XU225 offset[1] n202 NETTRAN_DUMMY_14768 NETTRAN_DUMMY_14769 CLKBUF_X1 
XU226 num_lzd_r[1] n203 NETTRAN_DUMMY_14770 NETTRAN_DUMMY_14771 INV_X1 
XU227 n203 n204 NETTRAN_DUMMY_14772 NETTRAN_DUMMY_14773 INV_X32 
XU228 n134 n205 NETTRAN_DUMMY_14774 NETTRAN_DUMMY_14775 BUF_X1 
XU229 offset[0] n206 NETTRAN_DUMMY_14776 NETTRAN_DUMMY_14777 INV_X32 
XU230 n206 n207 NETTRAN_DUMMY_14778 NETTRAN_DUMMY_14779 INV_X1 
XU231 n1098 n208 NETTRAN_DUMMY_14780 NETTRAN_DUMMY_14781 BUF_X1 
XU232 n1289 n209 NETTRAN_DUMMY_14782 NETTRAN_DUMMY_14783 BUF_X1 
XU233 n799 n210 NETTRAN_DUMMY_14784 NETTRAN_DUMMY_14785 BUF_X1 
XU234 c1_r1[17] n211 NETTRAN_DUMMY_14786 NETTRAN_DUMMY_14787 CLKBUF_X1 
XU235 n213 n212 NETTRAN_DUMMY_14788 NETTRAN_DUMMY_14789 CLKBUF_X1 
XU236 n211 n213 NETTRAN_DUMMY_14790 NETTRAN_DUMMY_14791 INV_X32 
XU237 n212 n214 NETTRAN_DUMMY_14792 NETTRAN_DUMMY_14793 INV_X32 
XU238 c1_r1[16] n215 NETTRAN_DUMMY_14794 NETTRAN_DUMMY_14795 CLKBUF_X1 
XU239 n217 n216 NETTRAN_DUMMY_14796 NETTRAN_DUMMY_14797 CLKBUF_X1 
XU240 n215 n217 NETTRAN_DUMMY_14798 NETTRAN_DUMMY_14799 INV_X32 
XU241 n216 n218 NETTRAN_DUMMY_14800 NETTRAN_DUMMY_14801 INV_X32 
XU242 c1_r1[15] n219 NETTRAN_DUMMY_14802 NETTRAN_DUMMY_14803 CLKBUF_X1 
XU243 n221 n220 NETTRAN_DUMMY_14804 NETTRAN_DUMMY_14805 CLKBUF_X1 
XU244 n219 n221 NETTRAN_DUMMY_14806 NETTRAN_DUMMY_14807 INV_X32 
XU245 n220 n222 NETTRAN_DUMMY_14808 NETTRAN_DUMMY_14809 INV_X32 
XU246 c1_r1[14] n223 NETTRAN_DUMMY_14810 NETTRAN_DUMMY_14811 CLKBUF_X1 
XU247 n225 n224 NETTRAN_DUMMY_14812 NETTRAN_DUMMY_14813 CLKBUF_X1 
XU248 n223 n225 NETTRAN_DUMMY_14814 NETTRAN_DUMMY_14815 INV_X32 
XU249 n224 n226 NETTRAN_DUMMY_14816 NETTRAN_DUMMY_14817 INV_X32 
XU250 c1_r1[13] n227 NETTRAN_DUMMY_14818 NETTRAN_DUMMY_14819 CLKBUF_X1 
XU251 n229 n228 NETTRAN_DUMMY_14820 NETTRAN_DUMMY_14821 CLKBUF_X1 
XU252 n227 n229 NETTRAN_DUMMY_14822 NETTRAN_DUMMY_14823 INV_X32 
XU253 n228 n230 NETTRAN_DUMMY_14824 NETTRAN_DUMMY_14825 INV_X32 
XU254 c1_r1[12] n231 NETTRAN_DUMMY_14826 NETTRAN_DUMMY_14827 CLKBUF_X1 
XU255 n233 n232 NETTRAN_DUMMY_14828 NETTRAN_DUMMY_14829 CLKBUF_X1 
XU256 n231 n233 NETTRAN_DUMMY_14830 NETTRAN_DUMMY_14831 INV_X32 
XU257 n232 n234 NETTRAN_DUMMY_14832 NETTRAN_DUMMY_14833 INV_X32 
XU258 c1_r1[11] n235 NETTRAN_DUMMY_14834 NETTRAN_DUMMY_14835 CLKBUF_X1 
XU259 n237 n236 NETTRAN_DUMMY_14836 NETTRAN_DUMMY_14837 CLKBUF_X1 
XU260 n235 n237 NETTRAN_DUMMY_14838 NETTRAN_DUMMY_14839 INV_X32 
XU261 n236 n238 NETTRAN_DUMMY_14840 NETTRAN_DUMMY_14841 INV_X32 
XU262 c1_r1[10] n239 NETTRAN_DUMMY_14842 NETTRAN_DUMMY_14843 CLKBUF_X1 
XU263 n241 n240 NETTRAN_DUMMY_14844 NETTRAN_DUMMY_14845 CLKBUF_X1 
XU264 n239 n241 NETTRAN_DUMMY_14846 NETTRAN_DUMMY_14847 INV_X32 
XU265 n240 n242 NETTRAN_DUMMY_14848 NETTRAN_DUMMY_14849 INV_X32 
XU266 c1_r1[9] n243 NETTRAN_DUMMY_14850 NETTRAN_DUMMY_14851 CLKBUF_X1 
XU267 n245 n244 NETTRAN_DUMMY_14852 NETTRAN_DUMMY_14853 CLKBUF_X1 
XU268 n243 n245 NETTRAN_DUMMY_14854 NETTRAN_DUMMY_14855 INV_X32 
XU269 n244 n246 NETTRAN_DUMMY_14856 NETTRAN_DUMMY_14857 INV_X32 
XU270 c1_r1[8] n247 NETTRAN_DUMMY_14858 NETTRAN_DUMMY_14859 CLKBUF_X1 
XU271 n249 n248 NETTRAN_DUMMY_14860 NETTRAN_DUMMY_14861 CLKBUF_X1 
XU272 n247 n249 NETTRAN_DUMMY_14862 NETTRAN_DUMMY_14863 INV_X32 
XU273 n248 n250 NETTRAN_DUMMY_14864 NETTRAN_DUMMY_14865 INV_X32 
XU274 c1_r1[7] n251 NETTRAN_DUMMY_14866 NETTRAN_DUMMY_14867 CLKBUF_X1 
XU275 n253 n252 NETTRAN_DUMMY_14868 NETTRAN_DUMMY_14869 CLKBUF_X1 
XU276 n251 n253 NETTRAN_DUMMY_14870 NETTRAN_DUMMY_14871 INV_X32 
XU277 n252 n254 NETTRAN_DUMMY_14872 NETTRAN_DUMMY_14873 INV_X32 
XU278 c1_r1[6] n255 NETTRAN_DUMMY_14874 NETTRAN_DUMMY_14875 CLKBUF_X1 
XU279 n257 n256 NETTRAN_DUMMY_14876 NETTRAN_DUMMY_14877 CLKBUF_X1 
XU280 n255 n257 NETTRAN_DUMMY_14878 NETTRAN_DUMMY_14879 INV_X32 
XU281 n256 n258 NETTRAN_DUMMY_14880 NETTRAN_DUMMY_14881 INV_X32 
XU282 c1_r1[5] n259 NETTRAN_DUMMY_14882 NETTRAN_DUMMY_14883 CLKBUF_X1 
XU283 n261 n260 NETTRAN_DUMMY_14884 NETTRAN_DUMMY_14885 CLKBUF_X1 
XU284 n259 n261 NETTRAN_DUMMY_14886 NETTRAN_DUMMY_14887 INV_X32 
XU285 n260 n262 NETTRAN_DUMMY_14888 NETTRAN_DUMMY_14889 INV_X32 
XU286 c1_r1[4] n263 NETTRAN_DUMMY_14890 NETTRAN_DUMMY_14891 CLKBUF_X1 
XU287 n265 n264 NETTRAN_DUMMY_14892 NETTRAN_DUMMY_14893 CLKBUF_X1 
XU288 n263 n265 NETTRAN_DUMMY_14894 NETTRAN_DUMMY_14895 INV_X32 
XU289 n264 n266 NETTRAN_DUMMY_14896 NETTRAN_DUMMY_14897 INV_X32 
XU290 c1_r1[3] n267 NETTRAN_DUMMY_14898 NETTRAN_DUMMY_14899 CLKBUF_X1 
XU291 n269 n268 NETTRAN_DUMMY_14900 NETTRAN_DUMMY_14901 CLKBUF_X1 
XU292 n267 n269 NETTRAN_DUMMY_14902 NETTRAN_DUMMY_14903 INV_X32 
XU293 n268 n270 NETTRAN_DUMMY_14904 NETTRAN_DUMMY_14905 INV_X32 
XU294 c1_r1[2] n271 NETTRAN_DUMMY_14906 NETTRAN_DUMMY_14907 CLKBUF_X1 
XU295 n150 n272 NETTRAN_DUMMY_14908 NETTRAN_DUMMY_14909 CLKBUF_X1 
XU296 n271 n273 NETTRAN_DUMMY_14910 NETTRAN_DUMMY_14911 INV_X32 
XU297 n272 n274 NETTRAN_DUMMY_14912 NETTRAN_DUMMY_14913 INV_X32 
XU298 c1_r1[1] n275 NETTRAN_DUMMY_14914 NETTRAN_DUMMY_14915 CLKBUF_X1 
XU299 n277 n276 NETTRAN_DUMMY_14916 NETTRAN_DUMMY_14917 CLKBUF_X1 
XU300 n275 n277 NETTRAN_DUMMY_14918 NETTRAN_DUMMY_14919 INV_X32 
XU301 n276 n278 NETTRAN_DUMMY_14920 NETTRAN_DUMMY_14921 INV_X32 
XU302 c1_r1[0] n279 NETTRAN_DUMMY_14922 NETTRAN_DUMMY_14923 CLKBUF_X1 
XU303 n281 n280 NETTRAN_DUMMY_14924 NETTRAN_DUMMY_14925 CLKBUF_X1 
XU304 n279 n281 NETTRAN_DUMMY_14926 NETTRAN_DUMMY_14927 INV_X32 
XU305 n280 n282 NETTRAN_DUMMY_14928 NETTRAN_DUMMY_14929 INV_X32 
XU306 x_r4[14] n283 NETTRAN_DUMMY_14930 NETTRAN_DUMMY_14931 CLKBUF_X1 
XU307 n285 n284 NETTRAN_DUMMY_14932 NETTRAN_DUMMY_14933 CLKBUF_X1 
XU308 n283 n285 NETTRAN_DUMMY_14934 NETTRAN_DUMMY_14935 INV_X32 
XU309 n284 n286 NETTRAN_DUMMY_14936 NETTRAN_DUMMY_14937 INV_X32 
XU310 x_r4[13] n287 NETTRAN_DUMMY_14938 NETTRAN_DUMMY_14939 CLKBUF_X1 
XU311 n289 n288 NETTRAN_DUMMY_14940 NETTRAN_DUMMY_14941 CLKBUF_X1 
XU312 n287 n289 NETTRAN_DUMMY_14942 NETTRAN_DUMMY_14943 INV_X32 
XU313 n288 n290 NETTRAN_DUMMY_14944 NETTRAN_DUMMY_14945 INV_X32 
XU314 x_r4[12] n291 NETTRAN_DUMMY_14946 NETTRAN_DUMMY_14947 CLKBUF_X1 
XU315 n293 n292 NETTRAN_DUMMY_14948 NETTRAN_DUMMY_14949 CLKBUF_X1 
XU316 n291 n293 NETTRAN_DUMMY_14950 NETTRAN_DUMMY_14951 INV_X32 
XU317 n292 n294 NETTRAN_DUMMY_14952 NETTRAN_DUMMY_14953 INV_X32 
XU318 x_r4[11] n295 NETTRAN_DUMMY_14954 NETTRAN_DUMMY_14955 CLKBUF_X1 
XU319 n297 n296 NETTRAN_DUMMY_14956 NETTRAN_DUMMY_14957 CLKBUF_X1 
XU320 n295 n297 NETTRAN_DUMMY_14958 NETTRAN_DUMMY_14959 INV_X32 
XU321 n296 n298 NETTRAN_DUMMY_14960 NETTRAN_DUMMY_14961 INV_X32 
XU322 x_r4[10] n299 NETTRAN_DUMMY_14962 NETTRAN_DUMMY_14963 CLKBUF_X1 
XU323 n301 n300 NETTRAN_DUMMY_14964 NETTRAN_DUMMY_14965 CLKBUF_X1 
XU324 n299 n301 NETTRAN_DUMMY_14966 NETTRAN_DUMMY_14967 INV_X32 
XU325 n300 n302 NETTRAN_DUMMY_14968 NETTRAN_DUMMY_14969 INV_X32 
XU326 x_r4[9] n303 NETTRAN_DUMMY_14970 NETTRAN_DUMMY_14971 CLKBUF_X1 
XU327 n305 n304 NETTRAN_DUMMY_14972 NETTRAN_DUMMY_14973 CLKBUF_X1 
XU328 n303 n305 NETTRAN_DUMMY_14974 NETTRAN_DUMMY_14975 INV_X32 
XU329 n304 n306 NETTRAN_DUMMY_14976 NETTRAN_DUMMY_14977 INV_X32 
XU330 x_r4[8] n307 NETTRAN_DUMMY_14978 NETTRAN_DUMMY_14979 CLKBUF_X1 
XU331 n309 n308 NETTRAN_DUMMY_14980 NETTRAN_DUMMY_14981 CLKBUF_X1 
XU332 n307 n309 NETTRAN_DUMMY_14982 NETTRAN_DUMMY_14983 INV_X32 
XU333 n308 n310 NETTRAN_DUMMY_14984 NETTRAN_DUMMY_14985 INV_X32 
XU334 x_r4[7] n311 NETTRAN_DUMMY_14986 NETTRAN_DUMMY_14987 CLKBUF_X1 
XU335 n313 n312 NETTRAN_DUMMY_14988 NETTRAN_DUMMY_14989 CLKBUF_X1 
XU336 n311 n313 NETTRAN_DUMMY_14990 NETTRAN_DUMMY_14991 INV_X32 
XU337 n312 n314 NETTRAN_DUMMY_14992 NETTRAN_DUMMY_14993 INV_X32 
XU338 x_r4[6] n315 NETTRAN_DUMMY_14994 NETTRAN_DUMMY_14995 CLKBUF_X1 
XU339 n317 n316 NETTRAN_DUMMY_14996 NETTRAN_DUMMY_14997 CLKBUF_X1 
XU340 n315 n317 NETTRAN_DUMMY_14998 NETTRAN_DUMMY_14999 INV_X32 
XU341 n316 n318 NETTRAN_DUMMY_15000 NETTRAN_DUMMY_15001 INV_X32 
XU342 x_r4[5] n319 NETTRAN_DUMMY_15002 NETTRAN_DUMMY_15003 CLKBUF_X1 
XU343 n321 n320 NETTRAN_DUMMY_15004 NETTRAN_DUMMY_15005 CLKBUF_X1 
XU344 n319 n321 NETTRAN_DUMMY_15006 NETTRAN_DUMMY_15007 INV_X32 
XU345 n320 n322 NETTRAN_DUMMY_15008 NETTRAN_DUMMY_15009 INV_X32 
XU346 x_r4[4] n323 NETTRAN_DUMMY_15010 NETTRAN_DUMMY_15011 CLKBUF_X1 
XU347 n325 n324 NETTRAN_DUMMY_15012 NETTRAN_DUMMY_15013 CLKBUF_X1 
XU348 n323 n325 NETTRAN_DUMMY_15014 NETTRAN_DUMMY_15015 INV_X32 
XU349 n324 n326 NETTRAN_DUMMY_15016 NETTRAN_DUMMY_15017 INV_X32 
XU350 x_r4[3] n327 NETTRAN_DUMMY_15018 NETTRAN_DUMMY_15019 CLKBUF_X1 
XU351 n329 n328 NETTRAN_DUMMY_15020 NETTRAN_DUMMY_15021 CLKBUF_X1 
XU352 n327 n329 NETTRAN_DUMMY_15022 NETTRAN_DUMMY_15023 INV_X32 
XU353 n328 n330 NETTRAN_DUMMY_15024 NETTRAN_DUMMY_15025 INV_X32 
XU354 x_r4[2] n331 NETTRAN_DUMMY_15026 NETTRAN_DUMMY_15027 CLKBUF_X1 
XU355 n333 n332 NETTRAN_DUMMY_15028 NETTRAN_DUMMY_15029 CLKBUF_X1 
XU356 n331 n333 NETTRAN_DUMMY_15030 NETTRAN_DUMMY_15031 INV_X32 
XU357 n332 n334 NETTRAN_DUMMY_15032 NETTRAN_DUMMY_15033 INV_X32 
XU358 x_r4[1] n335 NETTRAN_DUMMY_15034 NETTRAN_DUMMY_15035 CLKBUF_X1 
XU359 n337 n336 NETTRAN_DUMMY_15036 NETTRAN_DUMMY_15037 CLKBUF_X1 
XU360 n335 n337 NETTRAN_DUMMY_15038 NETTRAN_DUMMY_15039 INV_X32 
XU361 n336 n338 NETTRAN_DUMMY_15040 NETTRAN_DUMMY_15041 INV_X32 
XU362 x_r4[0] n339 NETTRAN_DUMMY_15042 NETTRAN_DUMMY_15043 CLKBUF_X1 
XU363 n341 n340 NETTRAN_DUMMY_15044 NETTRAN_DUMMY_15045 CLKBUF_X1 
XU364 n339 n341 NETTRAN_DUMMY_15046 NETTRAN_DUMMY_15047 INV_X32 
XU365 n340 n342 NETTRAN_DUMMY_15048 NETTRAN_DUMMY_15049 INV_X32 
XU366 n346 n343 NETTRAN_DUMMY_15050 NETTRAN_DUMMY_15051 CLKBUF_X1 
XU367 n343 n344 NETTRAN_DUMMY_15052 NETTRAN_DUMMY_15053 INV_X32 
XU368 n344 n345 NETTRAN_DUMMY_15054 NETTRAN_DUMMY_15055 INV_X1 
XU369 n22 n346 NETTRAN_DUMMY_15056 NETTRAN_DUMMY_15057 INV_X1 
XU370 n345 n347 NETTRAN_DUMMY_15058 NETTRAN_DUMMY_15059 INV_X32 
XU371 n349 n348 NETTRAN_DUMMY_15060 NETTRAN_DUMMY_15061 CLKBUF_X1 
XU372 n352 n349 NETTRAN_DUMMY_15062 NETTRAN_DUMMY_15063 INV_X1 
XU373 n348 n350 NETTRAN_DUMMY_15064 NETTRAN_DUMMY_15065 INV_X32 
XU374 n1 n351 NETTRAN_DUMMY_15066 NETTRAN_DUMMY_15067 INV_X1 
XU375 n351 n352 NETTRAN_DUMMY_15068 NETTRAN_DUMMY_15069 INV_X32 
XU376 n356 n353 NETTRAN_DUMMY_15070 NETTRAN_DUMMY_15071 CLKBUF_X1 
XU377 n353 n354 NETTRAN_DUMMY_15072 NETTRAN_DUMMY_15073 INV_X32 
XU378 n354 n355 NETTRAN_DUMMY_15074 NETTRAN_DUMMY_15075 INV_X1 
XU379 n940 n356 NETTRAN_DUMMY_15076 NETTRAN_DUMMY_15077 INV_X1 
XU380 n355 n357 NETTRAN_DUMMY_15078 NETTRAN_DUMMY_15079 INV_X32 
XU381 n361 n358 NETTRAN_DUMMY_15080 NETTRAN_DUMMY_15081 CLKBUF_X1 
XU382 n358 n359 NETTRAN_DUMMY_15082 NETTRAN_DUMMY_15083 INV_X32 
XU383 n359 n360 NETTRAN_DUMMY_15084 NETTRAN_DUMMY_15085 INV_X1 
XU384 n930 n361 NETTRAN_DUMMY_15086 NETTRAN_DUMMY_15087 INV_X1 
XU385 n360 n362 NETTRAN_DUMMY_15088 NETTRAN_DUMMY_15089 INV_X32 
XU386 n366 n363 NETTRAN_DUMMY_15090 NETTRAN_DUMMY_15091 CLKBUF_X1 
XU387 n363 n364 NETTRAN_DUMMY_15092 NETTRAN_DUMMY_15093 INV_X32 
XU388 n364 n365 NETTRAN_DUMMY_15094 NETTRAN_DUMMY_15095 INV_X1 
XU389 n920 n366 NETTRAN_DUMMY_15096 NETTRAN_DUMMY_15097 INV_X1 
XU390 n365 n367 NETTRAN_DUMMY_15098 NETTRAN_DUMMY_15099 INV_X32 
XU391 n371 n368 NETTRAN_DUMMY_15100 NETTRAN_DUMMY_15101 CLKBUF_X1 
XU392 n368 n369 NETTRAN_DUMMY_15102 NETTRAN_DUMMY_15103 INV_X32 
XU393 n369 n370 NETTRAN_DUMMY_15104 NETTRAN_DUMMY_15105 INV_X1 
XU394 n911 n371 NETTRAN_DUMMY_15106 NETTRAN_DUMMY_15107 INV_X1 
XU395 n370 n372 NETTRAN_DUMMY_15108 NETTRAN_DUMMY_15109 INV_X32 
XU396 n376 n373 NETTRAN_DUMMY_15110 NETTRAN_DUMMY_15111 CLKBUF_X1 
XU397 n373 n374 NETTRAN_DUMMY_15112 NETTRAN_DUMMY_15113 INV_X32 
XU398 n374 n375 NETTRAN_DUMMY_15114 NETTRAN_DUMMY_15115 INV_X1 
XU399 n9000 n376 NETTRAN_DUMMY_15116 NETTRAN_DUMMY_15117 INV_X1 
XU400 n375 n377 NETTRAN_DUMMY_15118 NETTRAN_DUMMY_15119 INV_X32 
XU401 n381 n378 NETTRAN_DUMMY_15120 NETTRAN_DUMMY_15121 CLKBUF_X1 
XU402 n378 n379 NETTRAN_DUMMY_15122 NETTRAN_DUMMY_15123 INV_X32 
XU403 n379 n380 NETTRAN_DUMMY_15124 NETTRAN_DUMMY_15125 INV_X1 
XU404 n890 n381 NETTRAN_DUMMY_15126 NETTRAN_DUMMY_15127 INV_X1 
XU405 n380 n382 NETTRAN_DUMMY_15128 NETTRAN_DUMMY_15129 INV_X32 
XU406 N147 n383 NETTRAN_DUMMY_15130 NETTRAN_DUMMY_15131 CLKBUF_X1 
XU407 n385 n384 NETTRAN_DUMMY_15132 NETTRAN_DUMMY_15133 CLKBUF_X1 
XU408 n383 n385 NETTRAN_DUMMY_15134 NETTRAN_DUMMY_15135 INV_X32 
XU409 n384 n386 NETTRAN_DUMMY_15136 NETTRAN_DUMMY_15137 INV_X32 
XU410 n388 n387 NETTRAN_DUMMY_15138 NETTRAN_DUMMY_15139 CLKBUF_X1 
XU411 n391 n388 NETTRAN_DUMMY_15140 NETTRAN_DUMMY_15141 INV_X1 
XU412 n387 n389 NETTRAN_DUMMY_15142 NETTRAN_DUMMY_15143 INV_X32 
XU413 N197 n390 NETTRAN_DUMMY_15144 NETTRAN_DUMMY_15145 INV_X1 
XU414 n390 n391 NETTRAN_DUMMY_15146 NETTRAN_DUMMY_15147 INV_X32 
XU415 n394 n392 NETTRAN_DUMMY_15148 NETTRAN_DUMMY_15149 INV_X32 
XU416 n392 n393 NETTRAN_DUMMY_15150 NETTRAN_DUMMY_15151 INV_X1 
XU417 n397 n394 NETTRAN_DUMMY_15152 NETTRAN_DUMMY_15153 INV_X1 
XU418 n393 n395 NETTRAN_DUMMY_15154 NETTRAN_DUMMY_15155 INV_X32 
XU419 N196 n396 NETTRAN_DUMMY_15156 NETTRAN_DUMMY_15157 INV_X1 
XU420 n396 n397 NETTRAN_DUMMY_15158 NETTRAN_DUMMY_15159 INV_X32 
XU421 n399 n398 NETTRAN_DUMMY_15160 NETTRAN_DUMMY_15161 CLKBUF_X1 
XU422 n402 n399 NETTRAN_DUMMY_15162 NETTRAN_DUMMY_15163 INV_X1 
XU423 n398 n400 NETTRAN_DUMMY_15164 NETTRAN_DUMMY_15165 INV_X32 
XU424 N195 n401 NETTRAN_DUMMY_15166 NETTRAN_DUMMY_15167 INV_X1 
XU425 n401 n402 NETTRAN_DUMMY_15168 NETTRAN_DUMMY_15169 INV_X32 
XU426 n405 n403 NETTRAN_DUMMY_15170 NETTRAN_DUMMY_15171 CLKBUF_X1 
XU427 n406 n404 NETTRAN_DUMMY_15172 NETTRAN_DUMMY_15173 INV_X32 
XU428 n404 n405 NETTRAN_DUMMY_15174 NETTRAN_DUMMY_15175 INV_X1 
XU429 N194 n406 NETTRAN_DUMMY_15176 NETTRAN_DUMMY_15177 INV_X1 
XU430 n403 n407 NETTRAN_DUMMY_15178 NETTRAN_DUMMY_15179 INV_X32 
XU431 n410 n408 NETTRAN_DUMMY_15180 NETTRAN_DUMMY_15181 CLKBUF_X1 
XU432 n412 n409 NETTRAN_DUMMY_15182 NETTRAN_DUMMY_15183 INV_X1 
XU433 n409 n410 NETTRAN_DUMMY_15184 NETTRAN_DUMMY_15185 INV_X32 
XU434 N193 n411 NETTRAN_DUMMY_15186 NETTRAN_DUMMY_15187 INV_X1 
XU435 n411 n412 NETTRAN_DUMMY_15188 NETTRAN_DUMMY_15189 INV_X32 
XU436 N192 n413 NETTRAN_DUMMY_15190 NETTRAN_DUMMY_15191 BUF_X16 
XU437 n417 n414 NETTRAN_DUMMY_15192 NETTRAN_DUMMY_15193 INV_X1 
XU438 n414 n415 NETTRAN_DUMMY_15194 NETTRAN_DUMMY_15195 INV_X32 
XU439 n413 n416 NETTRAN_DUMMY_15196 NETTRAN_DUMMY_15197 INV_X1 
XU440 n416 n417 NETTRAN_DUMMY_15198 NETTRAN_DUMMY_15199 INV_X32 
XU441 n419 n418 NETTRAN_DUMMY_15200 NETTRAN_DUMMY_15201 CLKBUF_X1 
XU442 n422 n419 NETTRAN_DUMMY_15202 NETTRAN_DUMMY_15203 INV_X1 
XU443 n418 n420 NETTRAN_DUMMY_15204 NETTRAN_DUMMY_15205 INV_X32 
XU444 N191 n421 NETTRAN_DUMMY_15206 NETTRAN_DUMMY_15207 INV_X1 
XU445 n421 n422 NETTRAN_DUMMY_15208 NETTRAN_DUMMY_15209 INV_X32 
XU446 n424 n423 NETTRAN_DUMMY_15210 NETTRAN_DUMMY_15211 CLKBUF_X1 
XU447 n427 n424 NETTRAN_DUMMY_15212 NETTRAN_DUMMY_15213 INV_X1 
XU448 n423 n425 NETTRAN_DUMMY_15214 NETTRAN_DUMMY_15215 INV_X32 
XU449 N190 n426 NETTRAN_DUMMY_15216 NETTRAN_DUMMY_15217 INV_X1 
XU450 n426 n427 NETTRAN_DUMMY_15218 NETTRAN_DUMMY_15219 INV_X32 
XU451 n430 n428 NETTRAN_DUMMY_15220 NETTRAN_DUMMY_15221 INV_X32 
XU452 n428 n429 NETTRAN_DUMMY_15222 NETTRAN_DUMMY_15223 INV_X1 
XU453 n433 n430 NETTRAN_DUMMY_15224 NETTRAN_DUMMY_15225 INV_X1 
XU454 n429 n431 NETTRAN_DUMMY_15226 NETTRAN_DUMMY_15227 INV_X32 
XU455 N189 n432 NETTRAN_DUMMY_15228 NETTRAN_DUMMY_15229 INV_X1 
XU456 n432 n433 NETTRAN_DUMMY_15230 NETTRAN_DUMMY_15231 INV_X32 
XU457 n436 n434 NETTRAN_DUMMY_15232 NETTRAN_DUMMY_15233 INV_X32 
XU458 n434 n435 NETTRAN_DUMMY_15234 NETTRAN_DUMMY_15235 INV_X1 
XU459 n439 n436 NETTRAN_DUMMY_15236 NETTRAN_DUMMY_15237 INV_X1 
XU460 n435 n437 NETTRAN_DUMMY_15238 NETTRAN_DUMMY_15239 INV_X32 
XU461 N188 n438 NETTRAN_DUMMY_15240 NETTRAN_DUMMY_15241 INV_X1 
XU462 n438 n439 NETTRAN_DUMMY_15242 NETTRAN_DUMMY_15243 INV_X32 
XU463 n442 n440 NETTRAN_DUMMY_15244 NETTRAN_DUMMY_15245 INV_X32 
XU464 n440 n441 NETTRAN_DUMMY_15246 NETTRAN_DUMMY_15247 INV_X1 
XU465 n445 n442 NETTRAN_DUMMY_15248 NETTRAN_DUMMY_15249 INV_X1 
XU466 n441 n443 NETTRAN_DUMMY_15250 NETTRAN_DUMMY_15251 INV_X32 
XU467 N187 n444 NETTRAN_DUMMY_15252 NETTRAN_DUMMY_15253 INV_X1 
XU468 n444 n445 NETTRAN_DUMMY_15254 NETTRAN_DUMMY_15255 INV_X32 
XU469 n448 n446 NETTRAN_DUMMY_15256 NETTRAN_DUMMY_15257 CLKBUF_X1 
XU470 n450 n447 NETTRAN_DUMMY_15258 NETTRAN_DUMMY_15259 INV_X1 
XU471 n447 n448 NETTRAN_DUMMY_15260 NETTRAN_DUMMY_15261 INV_X32 
XU472 N186 n449 NETTRAN_DUMMY_15262 NETTRAN_DUMMY_15263 INV_X1 
XU473 n449 n450 NETTRAN_DUMMY_15264 NETTRAN_DUMMY_15265 INV_X32 
XU474 n454 n451 NETTRAN_DUMMY_15266 NETTRAN_DUMMY_15267 INV_X1 
XU475 n451 n452 NETTRAN_DUMMY_15268 NETTRAN_DUMMY_15269 INV_X32 
XU476 N185 n453 NETTRAN_DUMMY_15270 NETTRAN_DUMMY_15271 INV_X1 
XU477 n453 n454 NETTRAN_DUMMY_15272 NETTRAN_DUMMY_15273 INV_X32 
XU478 n458 n455 NETTRAN_DUMMY_15274 NETTRAN_DUMMY_15275 INV_X1 
XU479 n455 n456 NETTRAN_DUMMY_15276 NETTRAN_DUMMY_15277 INV_X32 
XU480 n460 n457 NETTRAN_DUMMY_15278 NETTRAN_DUMMY_15279 INV_X1 
XU481 n457 n458 NETTRAN_DUMMY_15280 NETTRAN_DUMMY_15281 INV_X32 
XU482 N184 n459 NETTRAN_DUMMY_15282 NETTRAN_DUMMY_15283 INV_X1 
XU483 n459 n460 NETTRAN_DUMMY_15284 NETTRAN_DUMMY_15285 INV_X32 
XU484 n464 n461 NETTRAN_DUMMY_15286 NETTRAN_DUMMY_15287 INV_X1 
XU485 n461 n462 NETTRAN_DUMMY_15288 NETTRAN_DUMMY_15289 INV_X32 
XU486 n466 n463 NETTRAN_DUMMY_15290 NETTRAN_DUMMY_15291 INV_X1 
XU487 n463 n464 NETTRAN_DUMMY_15292 NETTRAN_DUMMY_15293 INV_X32 
XU488 N183 n465 NETTRAN_DUMMY_15294 NETTRAN_DUMMY_15295 INV_X1 
XU489 n465 n466 NETTRAN_DUMMY_15296 NETTRAN_DUMMY_15297 INV_X32 
XU490 n469 n467 NETTRAN_DUMMY_15298 NETTRAN_DUMMY_15299 INV_X32 
XU491 n467 n468 NETTRAN_DUMMY_15300 NETTRAN_DUMMY_15301 INV_X1 
XU492 n472 n469 NETTRAN_DUMMY_15302 NETTRAN_DUMMY_15303 INV_X1 
XU493 n468 n470 NETTRAN_DUMMY_15304 NETTRAN_DUMMY_15305 INV_X32 
XU494 N182 n471 NETTRAN_DUMMY_15306 NETTRAN_DUMMY_15307 INV_X1 
XU495 n471 n472 NETTRAN_DUMMY_15308 NETTRAN_DUMMY_15309 INV_X32 
XU496 c0_r2[8] n473 NETTRAN_DUMMY_15310 NETTRAN_DUMMY_15311 CLKBUF_X1 
XU497 n475 n474 NETTRAN_DUMMY_15312 NETTRAN_DUMMY_15313 CLKBUF_X1 
XU498 n473 n475 NETTRAN_DUMMY_15314 NETTRAN_DUMMY_15315 INV_X32 
XU499 n474 n476 NETTRAN_DUMMY_15316 NETTRAN_DUMMY_15317 INV_X32 
XU500 c0_r3[8] n477 NETTRAN_DUMMY_15318 NETTRAN_DUMMY_15319 CLKBUF_X1 
XU501 n479 n478 NETTRAN_DUMMY_15320 NETTRAN_DUMMY_15321 CLKBUF_X1 
XU502 n477 n479 NETTRAN_DUMMY_15322 NETTRAN_DUMMY_15323 INV_X32 
XU503 n478 n480 NETTRAN_DUMMY_15324 NETTRAN_DUMMY_15325 INV_X32 
XU504 c0_r1[7] n481 NETTRAN_DUMMY_15326 NETTRAN_DUMMY_15327 CLKBUF_X1 
XU505 n483 n482 NETTRAN_DUMMY_15328 NETTRAN_DUMMY_15329 CLKBUF_X1 
XU506 n481 n483 NETTRAN_DUMMY_15330 NETTRAN_DUMMY_15331 INV_X32 
XU507 n482 n484 NETTRAN_DUMMY_15332 NETTRAN_DUMMY_15333 INV_X32 
XU508 c0_r2[7] n485 NETTRAN_DUMMY_15334 NETTRAN_DUMMY_15335 CLKBUF_X1 
XU509 n487 n486 NETTRAN_DUMMY_15336 NETTRAN_DUMMY_15337 CLKBUF_X1 
XU510 n485 n487 NETTRAN_DUMMY_15338 NETTRAN_DUMMY_15339 INV_X32 
XU511 n486 n488 NETTRAN_DUMMY_15340 NETTRAN_DUMMY_15341 INV_X32 
XU512 c0_r3[7] n489 NETTRAN_DUMMY_15342 NETTRAN_DUMMY_15343 CLKBUF_X1 
XU513 n491 n490 NETTRAN_DUMMY_15344 NETTRAN_DUMMY_15345 CLKBUF_X1 
XU514 n489 n491 NETTRAN_DUMMY_15346 NETTRAN_DUMMY_15347 INV_X32 
XU515 n490 n492 NETTRAN_DUMMY_15348 NETTRAN_DUMMY_15349 INV_X32 
XU516 c0_r1[6] n493 NETTRAN_DUMMY_15350 NETTRAN_DUMMY_15351 CLKBUF_X1 
XU517 n495 n494 NETTRAN_DUMMY_15352 NETTRAN_DUMMY_15353 CLKBUF_X1 
XU518 n493 n495 NETTRAN_DUMMY_15354 NETTRAN_DUMMY_15355 INV_X32 
XU519 n494 n496 NETTRAN_DUMMY_15356 NETTRAN_DUMMY_15357 INV_X32 
XU520 c0_r2[6] n497 NETTRAN_DUMMY_15358 NETTRAN_DUMMY_15359 CLKBUF_X1 
XU521 n499 n498 NETTRAN_DUMMY_15360 NETTRAN_DUMMY_15361 CLKBUF_X1 
XU522 n497 n499 NETTRAN_DUMMY_15362 NETTRAN_DUMMY_15363 INV_X32 
XU523 n498 n500 NETTRAN_DUMMY_15364 NETTRAN_DUMMY_15365 INV_X32 
XU524 c0_r3[6] n501 NETTRAN_DUMMY_15366 NETTRAN_DUMMY_15367 CLKBUF_X1 
XU525 n503 n502 NETTRAN_DUMMY_15368 NETTRAN_DUMMY_15369 CLKBUF_X1 
XU526 n501 n503 NETTRAN_DUMMY_15370 NETTRAN_DUMMY_15371 INV_X32 
XU527 n502 n504 NETTRAN_DUMMY_15372 NETTRAN_DUMMY_15373 INV_X32 
XU528 c0_r1[5] n505 NETTRAN_DUMMY_15374 NETTRAN_DUMMY_15375 CLKBUF_X1 
XU529 n507 n506 NETTRAN_DUMMY_15376 NETTRAN_DUMMY_15377 CLKBUF_X1 
XU530 n505 n507 NETTRAN_DUMMY_15378 NETTRAN_DUMMY_15379 INV_X32 
XU531 n506 n508 NETTRAN_DUMMY_15380 NETTRAN_DUMMY_15381 INV_X32 
XU532 c0_r2[5] n509 NETTRAN_DUMMY_15382 NETTRAN_DUMMY_15383 CLKBUF_X1 
XU533 n511 n510 NETTRAN_DUMMY_15384 NETTRAN_DUMMY_15385 CLKBUF_X1 
XU534 n509 n511 NETTRAN_DUMMY_15386 NETTRAN_DUMMY_15387 INV_X32 
XU535 n510 n512 NETTRAN_DUMMY_15388 NETTRAN_DUMMY_15389 INV_X32 
XU536 c0_r3[5] n513 NETTRAN_DUMMY_15390 NETTRAN_DUMMY_15391 CLKBUF_X1 
XU537 n515 n514 NETTRAN_DUMMY_15392 NETTRAN_DUMMY_15393 CLKBUF_X1 
XU538 n513 n515 NETTRAN_DUMMY_15394 NETTRAN_DUMMY_15395 INV_X32 
XU539 n514 n516 NETTRAN_DUMMY_15396 NETTRAN_DUMMY_15397 INV_X32 
XU540 c0_r1[4] n517 NETTRAN_DUMMY_15398 NETTRAN_DUMMY_15399 CLKBUF_X1 
XU541 n519 n518 NETTRAN_DUMMY_15400 NETTRAN_DUMMY_15401 CLKBUF_X1 
XU542 n517 n519 NETTRAN_DUMMY_15402 NETTRAN_DUMMY_15403 INV_X32 
XU543 n518 n520 NETTRAN_DUMMY_15404 NETTRAN_DUMMY_15405 INV_X32 
XU544 c0_r2[4] n521 NETTRAN_DUMMY_15406 NETTRAN_DUMMY_15407 CLKBUF_X1 
XU545 n523 n522 NETTRAN_DUMMY_15408 NETTRAN_DUMMY_15409 CLKBUF_X1 
XU546 n521 n523 NETTRAN_DUMMY_15410 NETTRAN_DUMMY_15411 INV_X32 
XU547 n522 n524 NETTRAN_DUMMY_15412 NETTRAN_DUMMY_15413 INV_X32 
XU548 c0_r3[4] n525 NETTRAN_DUMMY_15414 NETTRAN_DUMMY_15415 CLKBUF_X1 
XU549 n527 n526 NETTRAN_DUMMY_15416 NETTRAN_DUMMY_15417 CLKBUF_X1 
XU550 n525 n527 NETTRAN_DUMMY_15418 NETTRAN_DUMMY_15419 INV_X32 
XU551 n526 n528 NETTRAN_DUMMY_15420 NETTRAN_DUMMY_15421 INV_X32 
XU552 c0_r1[3] n529 NETTRAN_DUMMY_15422 NETTRAN_DUMMY_15423 CLKBUF_X1 
XU553 n531 n530 NETTRAN_DUMMY_15424 NETTRAN_DUMMY_15425 CLKBUF_X1 
XU554 n529 n531 NETTRAN_DUMMY_15426 NETTRAN_DUMMY_15427 INV_X32 
XU555 n530 n532 NETTRAN_DUMMY_15428 NETTRAN_DUMMY_15429 INV_X32 
XU556 c0_r2[3] n533 NETTRAN_DUMMY_15430 NETTRAN_DUMMY_15431 CLKBUF_X1 
XU557 n535 n534 NETTRAN_DUMMY_15432 NETTRAN_DUMMY_15433 CLKBUF_X1 
XU558 n533 n535 NETTRAN_DUMMY_15434 NETTRAN_DUMMY_15435 INV_X32 
XU559 n534 n536 NETTRAN_DUMMY_15436 NETTRAN_DUMMY_15437 INV_X32 
XU560 c0_r3[3] n537 NETTRAN_DUMMY_15438 NETTRAN_DUMMY_15439 CLKBUF_X1 
XU561 n539 n538 NETTRAN_DUMMY_15440 NETTRAN_DUMMY_15441 CLKBUF_X1 
XU562 n537 n539 NETTRAN_DUMMY_15442 NETTRAN_DUMMY_15443 INV_X32 
XU563 n538 n540 NETTRAN_DUMMY_15444 NETTRAN_DUMMY_15445 INV_X32 
XU564 c0_r1[2] n541 NETTRAN_DUMMY_15446 NETTRAN_DUMMY_15447 CLKBUF_X1 
XU565 n543 n542 NETTRAN_DUMMY_15448 NETTRAN_DUMMY_15449 CLKBUF_X1 
XU566 n541 n543 NETTRAN_DUMMY_15450 NETTRAN_DUMMY_15451 INV_X32 
XU567 n542 n544 NETTRAN_DUMMY_15452 NETTRAN_DUMMY_15453 INV_X32 
XU568 c0_r2[2] n545 NETTRAN_DUMMY_15454 NETTRAN_DUMMY_15455 CLKBUF_X1 
XU569 n547 n546 NETTRAN_DUMMY_15456 NETTRAN_DUMMY_15457 CLKBUF_X1 
XU570 n545 n547 NETTRAN_DUMMY_15458 NETTRAN_DUMMY_15459 INV_X32 
XU571 n546 n548 NETTRAN_DUMMY_15460 NETTRAN_DUMMY_15461 INV_X32 
XU572 c0_r3[2] n549 NETTRAN_DUMMY_15462 NETTRAN_DUMMY_15463 CLKBUF_X1 
XU573 n551 n550 NETTRAN_DUMMY_15464 NETTRAN_DUMMY_15465 CLKBUF_X1 
XU574 n549 n551 NETTRAN_DUMMY_15466 NETTRAN_DUMMY_15467 INV_X32 
XU575 n550 n552 NETTRAN_DUMMY_15468 NETTRAN_DUMMY_15469 INV_X32 
XU576 c0_r1[1] n553 NETTRAN_DUMMY_15470 NETTRAN_DUMMY_15471 CLKBUF_X1 
XU577 n555 n554 NETTRAN_DUMMY_15472 NETTRAN_DUMMY_15473 CLKBUF_X1 
XU578 n553 n555 NETTRAN_DUMMY_15474 NETTRAN_DUMMY_15475 INV_X32 
XU579 n554 n556 NETTRAN_DUMMY_15476 NETTRAN_DUMMY_15477 INV_X32 
XU580 c0_r2[1] n557 NETTRAN_DUMMY_15478 NETTRAN_DUMMY_15479 CLKBUF_X1 
XU581 n559 n558 NETTRAN_DUMMY_15480 NETTRAN_DUMMY_15481 CLKBUF_X1 
XU582 n557 n559 NETTRAN_DUMMY_15482 NETTRAN_DUMMY_15483 INV_X32 
XU583 n558 n560 NETTRAN_DUMMY_15484 NETTRAN_DUMMY_15485 INV_X32 
XU584 c0_r3[1] n561 NETTRAN_DUMMY_15486 NETTRAN_DUMMY_15487 CLKBUF_X1 
XU585 n563 n562 NETTRAN_DUMMY_15488 NETTRAN_DUMMY_15489 CLKBUF_X1 
XU586 n561 n563 NETTRAN_DUMMY_15490 NETTRAN_DUMMY_15491 INV_X32 
XU587 n562 n564 NETTRAN_DUMMY_15492 NETTRAN_DUMMY_15493 INV_X32 
XU588 c0_r1[0] n565 NETTRAN_DUMMY_15494 NETTRAN_DUMMY_15495 CLKBUF_X1 
XU589 n567 n566 NETTRAN_DUMMY_15496 NETTRAN_DUMMY_15497 CLKBUF_X1 
XU590 n565 n567 NETTRAN_DUMMY_15498 NETTRAN_DUMMY_15499 INV_X32 
XU591 n566 n568 NETTRAN_DUMMY_15500 NETTRAN_DUMMY_15501 INV_X32 
XU592 c0_r2[0] n569 NETTRAN_DUMMY_15502 NETTRAN_DUMMY_15503 CLKBUF_X1 
XU593 n571 n570 NETTRAN_DUMMY_15504 NETTRAN_DUMMY_15505 CLKBUF_X1 
XU594 n569 n571 NETTRAN_DUMMY_15506 NETTRAN_DUMMY_15507 INV_X32 
XU595 n570 n572 NETTRAN_DUMMY_15508 NETTRAN_DUMMY_15509 INV_X32 
XU596 c0_r3[0] n573 NETTRAN_DUMMY_15510 NETTRAN_DUMMY_15511 CLKBUF_X1 
XU597 n575 n574 NETTRAN_DUMMY_15512 NETTRAN_DUMMY_15513 CLKBUF_X1 
XU598 n573 n575 NETTRAN_DUMMY_15514 NETTRAN_DUMMY_15515 INV_X32 
XU599 n574 n576 NETTRAN_DUMMY_15516 NETTRAN_DUMMY_15517 INV_X32 
XU600 c0_r4[17] n577 NETTRAN_DUMMY_15518 NETTRAN_DUMMY_15519 CLKBUF_X1 
XU601 n579 n578 NETTRAN_DUMMY_15520 NETTRAN_DUMMY_15521 CLKBUF_X1 
XU602 n577 n579 NETTRAN_DUMMY_15522 NETTRAN_DUMMY_15523 INV_X32 
XU603 n578 n580 NETTRAN_DUMMY_15524 NETTRAN_DUMMY_15525 INV_X32 
XU604 c0_r4[16] n581 NETTRAN_DUMMY_15526 NETTRAN_DUMMY_15527 CLKBUF_X1 
XU605 n583 n582 NETTRAN_DUMMY_15528 NETTRAN_DUMMY_15529 CLKBUF_X1 
XU606 n581 n583 NETTRAN_DUMMY_15530 NETTRAN_DUMMY_15531 INV_X32 
XU607 n582 n584 NETTRAN_DUMMY_15532 NETTRAN_DUMMY_15533 INV_X32 
XU608 c0_r4[15] n585 NETTRAN_DUMMY_15534 NETTRAN_DUMMY_15535 CLKBUF_X1 
XU609 n587 n586 NETTRAN_DUMMY_15536 NETTRAN_DUMMY_15537 CLKBUF_X1 
XU610 n585 n587 NETTRAN_DUMMY_15538 NETTRAN_DUMMY_15539 INV_X32 
XU611 n586 n588 NETTRAN_DUMMY_15540 NETTRAN_DUMMY_15541 INV_X32 
XU612 n592 n589 NETTRAN_DUMMY_15542 NETTRAN_DUMMY_15543 CLKBUF_X1 
XU613 n591 n590 NETTRAN_DUMMY_15544 NETTRAN_DUMMY_15545 CLKBUF_X1 
XU614 c0_r4[14] n591 NETTRAN_DUMMY_15546 NETTRAN_DUMMY_15547 INV_X32 
XU615 n590 n592 NETTRAN_DUMMY_15548 NETTRAN_DUMMY_15549 INV_X32 
XU616 c0_r4[13] n593 NETTRAN_DUMMY_15550 NETTRAN_DUMMY_15551 CLKBUF_X1 
XU617 n595 n594 NETTRAN_DUMMY_15552 NETTRAN_DUMMY_15553 CLKBUF_X1 
XU618 n593 n595 NETTRAN_DUMMY_15554 NETTRAN_DUMMY_15555 INV_X32 
XU619 n594 n596 NETTRAN_DUMMY_15556 NETTRAN_DUMMY_15557 INV_X32 
XU620 c0_r4[12] n597 NETTRAN_DUMMY_15558 NETTRAN_DUMMY_15559 CLKBUF_X1 
XU621 n599 n598 NETTRAN_DUMMY_15560 NETTRAN_DUMMY_15561 CLKBUF_X1 
XU622 n597 n599 NETTRAN_DUMMY_15562 NETTRAN_DUMMY_15563 INV_X32 
XU623 n598 n601 NETTRAN_DUMMY_15564 NETTRAN_DUMMY_15565 INV_X32 
XU624 c0_r4[11] n602 NETTRAN_DUMMY_15566 NETTRAN_DUMMY_15567 CLKBUF_X1 
XU625 n604 n603 NETTRAN_DUMMY_15568 NETTRAN_DUMMY_15569 CLKBUF_X1 
XU626 n602 n604 NETTRAN_DUMMY_15570 NETTRAN_DUMMY_15571 INV_X32 
XU627 n603 n605 NETTRAN_DUMMY_15572 NETTRAN_DUMMY_15573 INV_X32 
XU628 c0_r4[10] n606 NETTRAN_DUMMY_15574 NETTRAN_DUMMY_15575 CLKBUF_X1 
XU629 n608 n607 NETTRAN_DUMMY_15576 NETTRAN_DUMMY_15577 CLKBUF_X1 
XU630 n606 n608 NETTRAN_DUMMY_15578 NETTRAN_DUMMY_15579 INV_X32 
XU631 n607 n609 NETTRAN_DUMMY_15580 NETTRAN_DUMMY_15581 INV_X32 
XU632 c0_r4[9] n612 NETTRAN_DUMMY_15582 NETTRAN_DUMMY_15583 CLKBUF_X1 
XU633 n614 n613 NETTRAN_DUMMY_15584 NETTRAN_DUMMY_15585 CLKBUF_X1 
XU634 n612 n614 NETTRAN_DUMMY_15586 NETTRAN_DUMMY_15587 INV_X32 
XU635 n613 n615 NETTRAN_DUMMY_15588 NETTRAN_DUMMY_15589 INV_X32 
XU636 c0_r4[8] n616 NETTRAN_DUMMY_15590 NETTRAN_DUMMY_15591 CLKBUF_X1 
XU637 n618 n617 NETTRAN_DUMMY_15592 NETTRAN_DUMMY_15593 CLKBUF_X1 
XU638 n616 n618 NETTRAN_DUMMY_15594 NETTRAN_DUMMY_15595 INV_X32 
XU639 n617 n619 NETTRAN_DUMMY_15596 NETTRAN_DUMMY_15597 INV_X32 
XU640 c0_r4[7] n621 NETTRAN_DUMMY_15598 NETTRAN_DUMMY_15599 CLKBUF_X1 
XU641 n623 n622 NETTRAN_DUMMY_15600 NETTRAN_DUMMY_15601 CLKBUF_X1 
XU642 n621 n623 NETTRAN_DUMMY_15602 NETTRAN_DUMMY_15603 INV_X32 
XU643 n622 n624 NETTRAN_DUMMY_15604 NETTRAN_DUMMY_15605 INV_X32 
XU644 c0_r4[6] n625 NETTRAN_DUMMY_15606 NETTRAN_DUMMY_15607 CLKBUF_X1 
XU645 n627 n626 NETTRAN_DUMMY_15608 NETTRAN_DUMMY_15609 CLKBUF_X1 
XU646 n625 n627 NETTRAN_DUMMY_15610 NETTRAN_DUMMY_15611 INV_X32 
XU647 n626 n628 NETTRAN_DUMMY_15612 NETTRAN_DUMMY_15613 INV_X32 
XU648 c0_r4[5] n629 NETTRAN_DUMMY_15614 NETTRAN_DUMMY_15615 CLKBUF_X1 
XU649 n632 n631 NETTRAN_DUMMY_15616 NETTRAN_DUMMY_15617 CLKBUF_X1 
XU650 n629 n632 NETTRAN_DUMMY_15618 NETTRAN_DUMMY_15619 INV_X32 
XU651 n631 n633 NETTRAN_DUMMY_15620 NETTRAN_DUMMY_15621 INV_X32 
XU652 c0_r4[4] n634 NETTRAN_DUMMY_15622 NETTRAN_DUMMY_15623 CLKBUF_X1 
XU653 n636 n635 NETTRAN_DUMMY_15624 NETTRAN_DUMMY_15625 CLKBUF_X1 
XU654 n634 n636 NETTRAN_DUMMY_15626 NETTRAN_DUMMY_15627 INV_X32 
XU655 n635 n637 NETTRAN_DUMMY_15628 NETTRAN_DUMMY_15629 INV_X32 
XU656 c0_r4[3] n638 NETTRAN_DUMMY_15630 NETTRAN_DUMMY_15631 CLKBUF_X1 
XU657 n641 n639 NETTRAN_DUMMY_15632 NETTRAN_DUMMY_15633 CLKBUF_X1 
XU658 n638 n641 NETTRAN_DUMMY_15634 NETTRAN_DUMMY_15635 INV_X32 
XU659 n639 n642 NETTRAN_DUMMY_15636 NETTRAN_DUMMY_15637 INV_X32 
XU660 c0_r4[2] n643 NETTRAN_DUMMY_15638 NETTRAN_DUMMY_15639 CLKBUF_X1 
XU661 n645 n644 NETTRAN_DUMMY_15640 NETTRAN_DUMMY_15641 CLKBUF_X1 
XU662 n643 n645 NETTRAN_DUMMY_15642 NETTRAN_DUMMY_15643 INV_X32 
XU663 n644 n646 NETTRAN_DUMMY_15644 NETTRAN_DUMMY_15645 INV_X32 
XU664 c0_r4[1] n647 NETTRAN_DUMMY_15646 NETTRAN_DUMMY_15647 CLKBUF_X1 
XU665 n649 n648 NETTRAN_DUMMY_15648 NETTRAN_DUMMY_15649 CLKBUF_X1 
XU666 n647 n649 NETTRAN_DUMMY_15650 NETTRAN_DUMMY_15651 INV_X32 
XU667 n648 n651 NETTRAN_DUMMY_15652 NETTRAN_DUMMY_15653 INV_X32 
XU668 c0_r4[0] n652 NETTRAN_DUMMY_15654 NETTRAN_DUMMY_15655 CLKBUF_X1 
XU669 n654 n653 NETTRAN_DUMMY_15656 NETTRAN_DUMMY_15657 CLKBUF_X1 
XU670 n652 n654 NETTRAN_DUMMY_15658 NETTRAN_DUMMY_15659 INV_X32 
XU671 n653 n655 NETTRAN_DUMMY_15660 NETTRAN_DUMMY_15661 INV_X32 
XU672 sign_r[0] n656 NETTRAN_DUMMY_15662 NETTRAN_DUMMY_15663 CLKBUF_X1 
XU673 n658 n657 NETTRAN_DUMMY_15664 NETTRAN_DUMMY_15665 CLKBUF_X1 
XU674 n656 n658 NETTRAN_DUMMY_15666 NETTRAN_DUMMY_15667 INV_X32 
XU675 n657 n659 NETTRAN_DUMMY_15668 NETTRAN_DUMMY_15669 INV_X32 
XU676 sign_r[1] n661 NETTRAN_DUMMY_15670 NETTRAN_DUMMY_15671 CLKBUF_X1 
XU677 n663 n662 NETTRAN_DUMMY_15672 NETTRAN_DUMMY_15673 CLKBUF_X1 
XU678 n661 n663 NETTRAN_DUMMY_15674 NETTRAN_DUMMY_15675 INV_X32 
XU679 n662 n664 NETTRAN_DUMMY_15676 NETTRAN_DUMMY_15677 INV_X32 
XU680 sign_r[2] n665 NETTRAN_DUMMY_15678 NETTRAN_DUMMY_15679 CLKBUF_X1 
XU681 n667 n666 NETTRAN_DUMMY_15680 NETTRAN_DUMMY_15681 CLKBUF_X1 
XU682 n665 n667 NETTRAN_DUMMY_15682 NETTRAN_DUMMY_15683 INV_X32 
XU683 n666 n668 NETTRAN_DUMMY_15684 NETTRAN_DUMMY_15685 INV_X32 
XU684 sign_r[3] n669 NETTRAN_DUMMY_15686 NETTRAN_DUMMY_15687 CLKBUF_X1 
XU685 n672 n671 NETTRAN_DUMMY_15688 NETTRAN_DUMMY_15689 CLKBUF_X1 
XU686 n669 n672 NETTRAN_DUMMY_15690 NETTRAN_DUMMY_15691 INV_X32 
XU687 n671 n673 NETTRAN_DUMMY_15692 NETTRAN_DUMMY_15693 INV_X32 
XU688 sign_r[4] n674 NETTRAN_DUMMY_15694 NETTRAN_DUMMY_15695 CLKBUF_X1 
XU689 n676 n675 NETTRAN_DUMMY_15696 NETTRAN_DUMMY_15697 CLKBUF_X1 
XU690 n674 n676 NETTRAN_DUMMY_15698 NETTRAN_DUMMY_15699 INV_X32 
XU691 n675 n677 NETTRAN_DUMMY_15700 NETTRAN_DUMMY_15701 INV_X32 
XU692 n682 n678 NETTRAN_DUMMY_15702 NETTRAN_DUMMY_15703 BUF_X1 
XU693 n681 n679 NETTRAN_DUMMY_15704 NETTRAN_DUMMY_15705 CLKBUF_X1 
XU694 sign_r[5] n681 NETTRAN_DUMMY_15706 NETTRAN_DUMMY_15707 INV_X32 
XU695 n679 n682 NETTRAN_DUMMY_15708 NETTRAN_DUMMY_15709 INV_X32 
XU696 sign_r[6] n683 NETTRAN_DUMMY_15710 NETTRAN_DUMMY_15711 CLKBUF_X1 
XU697 n685 n684 NETTRAN_DUMMY_15712 NETTRAN_DUMMY_15713 CLKBUF_X1 
XU698 n683 n685 NETTRAN_DUMMY_15714 NETTRAN_DUMMY_15715 INV_X32 
XU699 n684 n686 NETTRAN_DUMMY_15716 NETTRAN_DUMMY_15717 INV_X32 
XU700 sign_r[7] n687 NETTRAN_DUMMY_15718 NETTRAN_DUMMY_15719 CLKBUF_X1 
XU701 n689 n688 NETTRAN_DUMMY_15720 NETTRAN_DUMMY_15721 CLKBUF_X1 
XU702 n687 n689 NETTRAN_DUMMY_15722 NETTRAN_DUMMY_15723 INV_X32 
XU703 n688 n691 NETTRAN_DUMMY_15724 NETTRAN_DUMMY_15725 INV_X32 
XU704 n695 n692 NETTRAN_DUMMY_15726 NETTRAN_DUMMY_15727 BUF_X1 
XU705 n694 n693 NETTRAN_DUMMY_15728 NETTRAN_DUMMY_15729 CLKBUF_X1 
XU706 N107 n694 NETTRAN_DUMMY_15730 NETTRAN_DUMMY_15731 INV_X32 
XU707 n693 n695 NETTRAN_DUMMY_15732 NETTRAN_DUMMY_15733 INV_X32 
XU708 N108 n696 NETTRAN_DUMMY_15734 NETTRAN_DUMMY_15735 CLKBUF_X1 
XU709 n698 n697 NETTRAN_DUMMY_15736 NETTRAN_DUMMY_15737 CLKBUF_X1 
XU710 n696 n698 NETTRAN_DUMMY_15738 NETTRAN_DUMMY_15739 INV_X32 
XU711 n697 n699 NETTRAN_DUMMY_15740 NETTRAN_DUMMY_15741 INV_X32 
XU712 valid_in_r[1] n701 NETTRAN_DUMMY_15742 NETTRAN_DUMMY_15743 CLKBUF_X1 
XU713 n703 n702 NETTRAN_DUMMY_15744 NETTRAN_DUMMY_15745 CLKBUF_X1 
XU714 n701 n703 NETTRAN_DUMMY_15746 NETTRAN_DUMMY_15747 INV_X32 
XU715 n702 n704 NETTRAN_DUMMY_15748 NETTRAN_DUMMY_15749 INV_X32 
XU716 N11010 n705 NETTRAN_DUMMY_15750 NETTRAN_DUMMY_15751 CLKBUF_X1 
XU717 n707 n706 NETTRAN_DUMMY_15752 NETTRAN_DUMMY_15753 CLKBUF_X1 
XU718 n705 n707 NETTRAN_DUMMY_15754 NETTRAN_DUMMY_15755 INV_X32 
XU719 n706 n708 NETTRAN_DUMMY_15756 NETTRAN_DUMMY_15757 INV_X32 
XU720 N111 n709 NETTRAN_DUMMY_15758 NETTRAN_DUMMY_15759 CLKBUF_X1 
XU721 n713 n712 NETTRAN_DUMMY_15760 NETTRAN_DUMMY_15761 CLKBUF_X1 
XU722 n709 n713 NETTRAN_DUMMY_15762 NETTRAN_DUMMY_15763 INV_X32 
XU723 n712 n714 NETTRAN_DUMMY_15764 NETTRAN_DUMMY_15765 INV_X32 
XU724 N112 n715 NETTRAN_DUMMY_15766 NETTRAN_DUMMY_15767 CLKBUF_X1 
XU725 n717 n716 NETTRAN_DUMMY_15768 NETTRAN_DUMMY_15769 CLKBUF_X1 
XU726 n715 n717 NETTRAN_DUMMY_15770 NETTRAN_DUMMY_15771 INV_X32 
XU727 n716 n718 NETTRAN_DUMMY_15772 NETTRAN_DUMMY_15773 INV_X32 
XU728 N113 n719 NETTRAN_DUMMY_15774 NETTRAN_DUMMY_15775 CLKBUF_X1 
XU729 n722 n721 NETTRAN_DUMMY_15776 NETTRAN_DUMMY_15777 CLKBUF_X1 
XU730 n719 n722 NETTRAN_DUMMY_15778 NETTRAN_DUMMY_15779 INV_X32 
XU731 n721 n723 NETTRAN_DUMMY_15780 NETTRAN_DUMMY_15781 INV_X32 
XU732 N114 n724 NETTRAN_DUMMY_15782 NETTRAN_DUMMY_15783 CLKBUF_X1 
XU733 n726 n725 NETTRAN_DUMMY_15784 NETTRAN_DUMMY_15785 CLKBUF_X1 
XU734 n724 n726 NETTRAN_DUMMY_15786 NETTRAN_DUMMY_15787 INV_X32 
XU735 n725 n727 NETTRAN_DUMMY_15788 NETTRAN_DUMMY_15789 INV_X32 
XU736 N115 n728 NETTRAN_DUMMY_15790 NETTRAN_DUMMY_15791 CLKBUF_X1 
XU737 n731 n729 NETTRAN_DUMMY_15792 NETTRAN_DUMMY_15793 CLKBUF_X1 
XU738 n728 n731 NETTRAN_DUMMY_15794 NETTRAN_DUMMY_15795 INV_X32 
XU739 n729 n732 NETTRAN_DUMMY_15796 NETTRAN_DUMMY_15797 INV_X32 
XU740 n736 n733 NETTRAN_DUMMY_15798 NETTRAN_DUMMY_15799 CLKBUF_X1 
XU741 n733 n734 NETTRAN_DUMMY_15800 NETTRAN_DUMMY_15801 INV_X32 
XU742 n734 n735 NETTRAN_DUMMY_15802 NETTRAN_DUMMY_15803 INV_X1 
XU743 n57 n736 NETTRAN_DUMMY_15804 NETTRAN_DUMMY_15805 INV_X1 
XU744 n735 n737 NETTRAN_DUMMY_15806 NETTRAN_DUMMY_15807 INV_X32 
XU745 n741 n738 NETTRAN_DUMMY_15808 NETTRAN_DUMMY_15809 CLKBUF_X1 
XU746 n742 n739 NETTRAN_DUMMY_15810 NETTRAN_DUMMY_15811 INV_X32 
XU747 n739 n741 NETTRAN_DUMMY_15812 NETTRAN_DUMMY_15813 INV_X1 
XU748 n28 n742 NETTRAN_DUMMY_15814 NETTRAN_DUMMY_15815 INV_X1 
XU749 n738 n743 NETTRAN_DUMMY_15816 NETTRAN_DUMMY_15817 INV_X32 
XU750 n746 n744 NETTRAN_DUMMY_15818 NETTRAN_DUMMY_15819 CLKBUF_X1 
XU751 n747 n745 NETTRAN_DUMMY_15820 NETTRAN_DUMMY_15821 INV_X32 
XU752 n745 n746 NETTRAN_DUMMY_15822 NETTRAN_DUMMY_15823 INV_X1 
XU753 n27 n747 NETTRAN_DUMMY_15824 NETTRAN_DUMMY_15825 INV_X1 
XU754 n744 n748 NETTRAN_DUMMY_15826 NETTRAN_DUMMY_15827 INV_X32 
XU755 n752 n749 NETTRAN_DUMMY_15828 NETTRAN_DUMMY_15829 CLKBUF_X1 
XU756 n753 n751 NETTRAN_DUMMY_15830 NETTRAN_DUMMY_15831 INV_X32 
XU757 n751 n752 NETTRAN_DUMMY_15832 NETTRAN_DUMMY_15833 INV_X1 
XU758 n26 n753 NETTRAN_DUMMY_15834 NETTRAN_DUMMY_15835 INV_X1 
XU759 n749 n754 NETTRAN_DUMMY_15836 NETTRAN_DUMMY_15837 INV_X32 
XU760 n759 n755 NETTRAN_DUMMY_15838 NETTRAN_DUMMY_15839 BUF_X1 
XU761 n758 n756 NETTRAN_DUMMY_15840 NETTRAN_DUMMY_15841 INV_X32 
XU762 n756 n757 NETTRAN_DUMMY_15842 NETTRAN_DUMMY_15843 INV_X1 
XU763 n25 n758 NETTRAN_DUMMY_15844 NETTRAN_DUMMY_15845 INV_X1 
XU764 n757 n759 NETTRAN_DUMMY_15846 NETTRAN_DUMMY_15847 INV_X32 
XU765 n764 n761 NETTRAN_DUMMY_15848 NETTRAN_DUMMY_15849 CLKBUF_X1 
XU766 n761 n762 NETTRAN_DUMMY_15850 NETTRAN_DUMMY_15851 INV_X32 
XU767 n762 n763 NETTRAN_DUMMY_15852 NETTRAN_DUMMY_15853 INV_X1 
XU768 n24 n764 NETTRAN_DUMMY_15854 NETTRAN_DUMMY_15855 INV_X1 
XU769 n763 n765 NETTRAN_DUMMY_15856 NETTRAN_DUMMY_15857 INV_X32 
XU770 n769 n766 NETTRAN_DUMMY_15858 NETTRAN_DUMMY_15859 CLKBUF_X1 
XU771 n766 n767 NETTRAN_DUMMY_15860 NETTRAN_DUMMY_15861 INV_X32 
XU772 n767 n768 NETTRAN_DUMMY_15862 NETTRAN_DUMMY_15863 INV_X1 
XU773 n23 n769 NETTRAN_DUMMY_15864 NETTRAN_DUMMY_15865 INV_X1 
XU774 n768 n771 NETTRAN_DUMMY_15866 NETTRAN_DUMMY_15867 INV_X32 
XU775 x_r2[7] n772 NETTRAN_DUMMY_15868 NETTRAN_DUMMY_15869 CLKBUF_X1 
XU776 n774 n773 NETTRAN_DUMMY_15870 NETTRAN_DUMMY_15871 CLKBUF_X1 
XU777 n772 n774 NETTRAN_DUMMY_15872 NETTRAN_DUMMY_15873 INV_X32 
XU778 n773 n775 NETTRAN_DUMMY_15874 NETTRAN_DUMMY_15875 INV_X32 
XU779 n777 n776 NETTRAN_DUMMY_15876 NETTRAN_DUMMY_15877 CLKBUF_X1 
XU780 n781 n777 NETTRAN_DUMMY_15878 NETTRAN_DUMMY_15879 INV_X1 
XU781 n776 n778 NETTRAN_DUMMY_15880 NETTRAN_DUMMY_15881 INV_X32 
XU782 N100 n779 NETTRAN_DUMMY_15882 NETTRAN_DUMMY_15883 INV_X1 
XU783 n779 n781 NETTRAN_DUMMY_15884 NETTRAN_DUMMY_15885 INV_X32 
XU784 x_r1[6] n782 NETTRAN_DUMMY_15886 NETTRAN_DUMMY_15887 CLKBUF_X1 
XU785 n784 n783 NETTRAN_DUMMY_15888 NETTRAN_DUMMY_15889 CLKBUF_X1 
XU786 n782 n784 NETTRAN_DUMMY_15890 NETTRAN_DUMMY_15891 INV_X32 
XU787 n783 n785 NETTRAN_DUMMY_15892 NETTRAN_DUMMY_15893 INV_X32 
XU788 x_r2[6] n786 NETTRAN_DUMMY_15894 NETTRAN_DUMMY_15895 CLKBUF_X1 
XU789 n788 n787 NETTRAN_DUMMY_15896 NETTRAN_DUMMY_15897 CLKBUF_X1 
XU790 n786 n788 NETTRAN_DUMMY_15898 NETTRAN_DUMMY_15899 INV_X32 
XU791 n787 n789 NETTRAN_DUMMY_15900 NETTRAN_DUMMY_15901 INV_X32 
XU792 n794 n791 NETTRAN_DUMMY_15902 NETTRAN_DUMMY_15903 CLKBUF_X1 
XU793 N101 n792 NETTRAN_DUMMY_15904 NETTRAN_DUMMY_15905 INV_X1 
XU794 n792 n793 NETTRAN_DUMMY_15906 NETTRAN_DUMMY_15907 INV_X32 
XU795 n793 n794 NETTRAN_DUMMY_15908 NETTRAN_DUMMY_15909 INV_X1 
XU796 n791 n795 NETTRAN_DUMMY_15910 NETTRAN_DUMMY_15911 INV_X32 
XU797 x_r1[5] n796 NETTRAN_DUMMY_15912 NETTRAN_DUMMY_15913 CLKBUF_X1 
XU798 n798 n797 NETTRAN_DUMMY_15914 NETTRAN_DUMMY_15915 CLKBUF_X1 
XU799 n796 n798 NETTRAN_DUMMY_15916 NETTRAN_DUMMY_15917 INV_X32 
XU800 n797 n799 NETTRAN_DUMMY_15918 NETTRAN_DUMMY_15919 INV_X32 
XU801 x_r2[5] n801 NETTRAN_DUMMY_15920 NETTRAN_DUMMY_15921 CLKBUF_X1 
XU802 n803 n802 NETTRAN_DUMMY_15922 NETTRAN_DUMMY_15923 CLKBUF_X1 
XU803 n801 n803 NETTRAN_DUMMY_15924 NETTRAN_DUMMY_15925 INV_X32 
XU804 n802 n804 NETTRAN_DUMMY_15926 NETTRAN_DUMMY_15927 INV_X32 
XU805 n806 n805 NETTRAN_DUMMY_15928 NETTRAN_DUMMY_15929 CLKBUF_X1 
XU806 N102 n806 NETTRAN_DUMMY_15930 NETTRAN_DUMMY_15931 INV_X1 
XU807 n805 n807 NETTRAN_DUMMY_15932 NETTRAN_DUMMY_15933 INV_X32 
XU808 n807 n808 NETTRAN_DUMMY_15934 NETTRAN_DUMMY_15935 INV_X1 
XU809 n808 n809 NETTRAN_DUMMY_15936 NETTRAN_DUMMY_15937 INV_X32 
XU810 x_r1[4] n812 NETTRAN_DUMMY_15938 NETTRAN_DUMMY_15939 CLKBUF_X1 
XU811 n814 n813 NETTRAN_DUMMY_15940 NETTRAN_DUMMY_15941 CLKBUF_X1 
XU812 n812 n814 NETTRAN_DUMMY_15942 NETTRAN_DUMMY_15943 INV_X32 
XU813 n813 n815 NETTRAN_DUMMY_15944 NETTRAN_DUMMY_15945 INV_X32 
XU814 x_r2[4] n816 NETTRAN_DUMMY_15946 NETTRAN_DUMMY_15947 CLKBUF_X1 
XU815 n818 n817 NETTRAN_DUMMY_15948 NETTRAN_DUMMY_15949 CLKBUF_X1 
XU816 n816 n818 NETTRAN_DUMMY_15950 NETTRAN_DUMMY_15951 INV_X32 
XU817 n817 n819 NETTRAN_DUMMY_15952 NETTRAN_DUMMY_15953 INV_X32 
XU818 n824 n821 NETTRAN_DUMMY_15954 NETTRAN_DUMMY_15955 CLKBUF_X1 
XU819 N103 n822 NETTRAN_DUMMY_15956 NETTRAN_DUMMY_15957 INV_X1 
XU820 n822 n823 NETTRAN_DUMMY_15958 NETTRAN_DUMMY_15959 INV_X32 
XU821 n823 n824 NETTRAN_DUMMY_15960 NETTRAN_DUMMY_15961 INV_X1 
XU822 n821 n825 NETTRAN_DUMMY_15962 NETTRAN_DUMMY_15963 INV_X32 
XU823 x_r1[3] n826 NETTRAN_DUMMY_15964 NETTRAN_DUMMY_15965 CLKBUF_X1 
XU824 n828 n827 NETTRAN_DUMMY_15966 NETTRAN_DUMMY_15967 CLKBUF_X1 
XU825 n826 n828 NETTRAN_DUMMY_15968 NETTRAN_DUMMY_15969 INV_X32 
XU826 n827 n829 NETTRAN_DUMMY_15970 NETTRAN_DUMMY_15971 INV_X32 
XU827 x_r2[3] n831 NETTRAN_DUMMY_15972 NETTRAN_DUMMY_15973 CLKBUF_X1 
XU828 n833 n832 NETTRAN_DUMMY_15974 NETTRAN_DUMMY_15975 CLKBUF_X1 
XU829 n831 n833 NETTRAN_DUMMY_15976 NETTRAN_DUMMY_15977 INV_X32 
XU830 n832 n834 NETTRAN_DUMMY_15978 NETTRAN_DUMMY_15979 INV_X32 
XU831 n837 n835 NETTRAN_DUMMY_15980 NETTRAN_DUMMY_15981 INV_X32 
XU832 n835 n836 NETTRAN_DUMMY_15982 NETTRAN_DUMMY_15983 INV_X1 
XU833 n841 n837 NETTRAN_DUMMY_15984 NETTRAN_DUMMY_15985 INV_X1 
XU834 n836 n838 NETTRAN_DUMMY_15986 NETTRAN_DUMMY_15987 INV_X32 
XU835 N104 n839 NETTRAN_DUMMY_15988 NETTRAN_DUMMY_15989 INV_X1 
XU836 n839 n841 NETTRAN_DUMMY_15990 NETTRAN_DUMMY_15991 INV_X32 
XU837 x_r1[2] n842 NETTRAN_DUMMY_15992 NETTRAN_DUMMY_15993 CLKBUF_X1 
XU838 n844 n843 NETTRAN_DUMMY_15994 NETTRAN_DUMMY_15995 CLKBUF_X1 
XU839 n842 n844 NETTRAN_DUMMY_15996 NETTRAN_DUMMY_15997 INV_X32 
XU840 n843 n845 NETTRAN_DUMMY_15998 NETTRAN_DUMMY_15999 INV_X32 
XU841 x_r2[2] n846 NETTRAN_DUMMY_16000 NETTRAN_DUMMY_16001 CLKBUF_X1 
XU842 n848 n847 NETTRAN_DUMMY_16002 NETTRAN_DUMMY_16003 CLKBUF_X1 
XU843 n846 n848 NETTRAN_DUMMY_16004 NETTRAN_DUMMY_16005 INV_X32 
XU844 n847 n849 NETTRAN_DUMMY_16006 NETTRAN_DUMMY_16007 INV_X32 
XU845 n854 n851 NETTRAN_DUMMY_16008 NETTRAN_DUMMY_16009 CLKBUF_X1 
XU846 N105 n852 NETTRAN_DUMMY_16010 NETTRAN_DUMMY_16011 INV_X1 
XU847 n852 n853 NETTRAN_DUMMY_16012 NETTRAN_DUMMY_16013 INV_X32 
XU848 n853 n854 NETTRAN_DUMMY_16014 NETTRAN_DUMMY_16015 INV_X1 
XU849 n851 n855 NETTRAN_DUMMY_16016 NETTRAN_DUMMY_16017 INV_X32 
XU850 x_r1[1] n856 NETTRAN_DUMMY_16018 NETTRAN_DUMMY_16019 CLKBUF_X1 
XU851 n858 n857 NETTRAN_DUMMY_16020 NETTRAN_DUMMY_16021 CLKBUF_X1 
XU852 n856 n858 NETTRAN_DUMMY_16022 NETTRAN_DUMMY_16023 INV_X32 
XU853 n857 n859 NETTRAN_DUMMY_16024 NETTRAN_DUMMY_16025 INV_X32 
XU854 x_r2[1] n861 NETTRAN_DUMMY_16026 NETTRAN_DUMMY_16027 CLKBUF_X1 
XU855 n863 n862 NETTRAN_DUMMY_16028 NETTRAN_DUMMY_16029 CLKBUF_X1 
XU856 n861 n863 NETTRAN_DUMMY_16030 NETTRAN_DUMMY_16031 INV_X32 
XU857 n862 n864 NETTRAN_DUMMY_16032 NETTRAN_DUMMY_16033 INV_X32 
XU858 n868 n865 NETTRAN_DUMMY_16034 NETTRAN_DUMMY_16035 INV_X1 
XU859 n865 n866 NETTRAN_DUMMY_16036 NETTRAN_DUMMY_16037 INV_X32 
XU860 n871 n867 NETTRAN_DUMMY_16038 NETTRAN_DUMMY_16039 INV_X1 
XU861 n867 n868 NETTRAN_DUMMY_16040 NETTRAN_DUMMY_16041 INV_X32 
XU862 N106 n869 NETTRAN_DUMMY_16042 NETTRAN_DUMMY_16043 INV_X1 
XU863 n869 n871 NETTRAN_DUMMY_16044 NETTRAN_DUMMY_16045 INV_X32 
XU864 x_r1[0] n872 NETTRAN_DUMMY_16046 NETTRAN_DUMMY_16047 CLKBUF_X1 
XU865 n874 n873 NETTRAN_DUMMY_16048 NETTRAN_DUMMY_16049 CLKBUF_X1 
XU866 n872 n874 NETTRAN_DUMMY_16050 NETTRAN_DUMMY_16051 INV_X32 
XU867 n873 n875 NETTRAN_DUMMY_16052 NETTRAN_DUMMY_16053 INV_X32 
XU868 x_r2[0] n876 NETTRAN_DUMMY_16054 NETTRAN_DUMMY_16055 CLKBUF_X1 
XU869 n878 n877 NETTRAN_DUMMY_16056 NETTRAN_DUMMY_16057 CLKBUF_X1 
XU870 n876 n878 NETTRAN_DUMMY_16058 NETTRAN_DUMMY_16059 INV_X32 
XU871 n877 n879 NETTRAN_DUMMY_16060 NETTRAN_DUMMY_16061 INV_X32 
XU872 x_r3[14] n881 NETTRAN_DUMMY_16062 NETTRAN_DUMMY_16063 CLKBUF_X1 
XU873 n883 n882 NETTRAN_DUMMY_16064 NETTRAN_DUMMY_16065 CLKBUF_X1 
XU874 n881 n883 NETTRAN_DUMMY_16066 NETTRAN_DUMMY_16067 INV_X32 
XU875 n882 n884 NETTRAN_DUMMY_16068 NETTRAN_DUMMY_16069 INV_X32 
XU876 x_r3[13] n885 NETTRAN_DUMMY_16070 NETTRAN_DUMMY_16071 CLKBUF_X1 
XU877 n887 n886 NETTRAN_DUMMY_16072 NETTRAN_DUMMY_16073 CLKBUF_X1 
XU878 n885 n887 NETTRAN_DUMMY_16074 NETTRAN_DUMMY_16075 INV_X32 
XU879 n886 n888 NETTRAN_DUMMY_16076 NETTRAN_DUMMY_16077 INV_X32 
XU880 x_r3[12] n889 NETTRAN_DUMMY_16078 NETTRAN_DUMMY_16079 CLKBUF_X1 
XU881 n892 n891 NETTRAN_DUMMY_16080 NETTRAN_DUMMY_16081 CLKBUF_X1 
XU882 n889 n892 NETTRAN_DUMMY_16082 NETTRAN_DUMMY_16083 INV_X32 
XU883 n891 n893 NETTRAN_DUMMY_16084 NETTRAN_DUMMY_16085 INV_X32 
XU884 x_r3[11] n894 NETTRAN_DUMMY_16086 NETTRAN_DUMMY_16087 CLKBUF_X1 
XU885 n896 n895 NETTRAN_DUMMY_16088 NETTRAN_DUMMY_16089 CLKBUF_X1 
XU886 n894 n896 NETTRAN_DUMMY_16090 NETTRAN_DUMMY_16091 INV_X32 
XU887 n895 n897 NETTRAN_DUMMY_16092 NETTRAN_DUMMY_16093 INV_X32 
XU888 x_r3[10] n898 NETTRAN_DUMMY_16094 NETTRAN_DUMMY_16095 CLKBUF_X1 
XU889 n901 n899 NETTRAN_DUMMY_16096 NETTRAN_DUMMY_16097 CLKBUF_X1 
XU890 n898 n901 NETTRAN_DUMMY_16098 NETTRAN_DUMMY_16099 INV_X32 
XU891 n899 n902 NETTRAN_DUMMY_16100 NETTRAN_DUMMY_16101 INV_X32 
XU892 x_r3[9] n903 NETTRAN_DUMMY_16102 NETTRAN_DUMMY_16103 CLKBUF_X1 
XU893 n905 n904 NETTRAN_DUMMY_16104 NETTRAN_DUMMY_16105 CLKBUF_X1 
XU894 n903 n905 NETTRAN_DUMMY_16106 NETTRAN_DUMMY_16107 INV_X32 
XU895 n904 n906 NETTRAN_DUMMY_16108 NETTRAN_DUMMY_16109 INV_X32 
XU896 x_r3[8] n907 NETTRAN_DUMMY_16110 NETTRAN_DUMMY_16111 CLKBUF_X1 
XU897 n909 n908 NETTRAN_DUMMY_16112 NETTRAN_DUMMY_16113 CLKBUF_X1 
XU898 n907 n909 NETTRAN_DUMMY_16114 NETTRAN_DUMMY_16115 INV_X32 
XU899 n908 n912 NETTRAN_DUMMY_16116 NETTRAN_DUMMY_16117 INV_X32 
XU900 x_r3[7] n913 NETTRAN_DUMMY_16118 NETTRAN_DUMMY_16119 CLKBUF_X1 
XU901 n915 n914 NETTRAN_DUMMY_16120 NETTRAN_DUMMY_16121 CLKBUF_X1 
XU902 n913 n915 NETTRAN_DUMMY_16122 NETTRAN_DUMMY_16123 INV_X32 
XU903 n914 n916 NETTRAN_DUMMY_16124 NETTRAN_DUMMY_16125 INV_X32 
XU904 x_r3[6] n917 NETTRAN_DUMMY_16126 NETTRAN_DUMMY_16127 CLKBUF_X1 
XU905 n919 n918 NETTRAN_DUMMY_16128 NETTRAN_DUMMY_16129 CLKBUF_X1 
XU906 n917 n919 NETTRAN_DUMMY_16130 NETTRAN_DUMMY_16131 INV_X32 
XU907 n918 n921 NETTRAN_DUMMY_16132 NETTRAN_DUMMY_16133 INV_X32 
XU908 x_r3[5] n922 NETTRAN_DUMMY_16134 NETTRAN_DUMMY_16135 CLKBUF_X1 
XU909 n924 n923 NETTRAN_DUMMY_16136 NETTRAN_DUMMY_16137 CLKBUF_X1 
XU910 n922 n924 NETTRAN_DUMMY_16138 NETTRAN_DUMMY_16139 INV_X32 
XU911 n923 n925 NETTRAN_DUMMY_16140 NETTRAN_DUMMY_16141 INV_X32 
XU912 x_r3[4] n926 NETTRAN_DUMMY_16142 NETTRAN_DUMMY_16143 CLKBUF_X1 
XU913 n928 n927 NETTRAN_DUMMY_16144 NETTRAN_DUMMY_16145 CLKBUF_X1 
XU914 n926 n928 NETTRAN_DUMMY_16146 NETTRAN_DUMMY_16147 INV_X32 
XU915 n927 n929 NETTRAN_DUMMY_16148 NETTRAN_DUMMY_16149 INV_X32 
XU916 x_r3[3] n931 NETTRAN_DUMMY_16150 NETTRAN_DUMMY_16151 CLKBUF_X1 
XU917 n933 n932 NETTRAN_DUMMY_16152 NETTRAN_DUMMY_16153 CLKBUF_X1 
XU918 n931 n933 NETTRAN_DUMMY_16154 NETTRAN_DUMMY_16155 INV_X32 
XU919 n932 n934 NETTRAN_DUMMY_16156 NETTRAN_DUMMY_16157 INV_X32 
XU920 x_r3[2] n935 NETTRAN_DUMMY_16158 NETTRAN_DUMMY_16159 CLKBUF_X1 
XU921 n937 n936 NETTRAN_DUMMY_16160 NETTRAN_DUMMY_16161 CLKBUF_X1 
XU922 n935 n937 NETTRAN_DUMMY_16162 NETTRAN_DUMMY_16163 INV_X32 
XU923 n936 n938 NETTRAN_DUMMY_16164 NETTRAN_DUMMY_16165 INV_X32 
XU924 x_r3[1] n939 NETTRAN_DUMMY_16166 NETTRAN_DUMMY_16167 CLKBUF_X1 
XU925 n942 n941 NETTRAN_DUMMY_16168 NETTRAN_DUMMY_16169 CLKBUF_X1 
XU926 n939 n942 NETTRAN_DUMMY_16170 NETTRAN_DUMMY_16171 INV_X32 
XU927 n941 n943 NETTRAN_DUMMY_16172 NETTRAN_DUMMY_16173 INV_X32 
XU928 x_r3[0] n944 NETTRAN_DUMMY_16174 NETTRAN_DUMMY_16175 CLKBUF_X1 
XU929 n946 n945 NETTRAN_DUMMY_16176 NETTRAN_DUMMY_16177 CLKBUF_X1 
XU930 n944 n946 NETTRAN_DUMMY_16178 NETTRAN_DUMMY_16179 INV_X32 
XU931 n945 n947 NETTRAN_DUMMY_16180 NETTRAN_DUMMY_16181 INV_X32 
XU932 c0_r1[17] n948 NETTRAN_DUMMY_16182 NETTRAN_DUMMY_16183 CLKBUF_X1 
XU933 n951 n949 NETTRAN_DUMMY_16184 NETTRAN_DUMMY_16185 CLKBUF_X1 
XU934 n948 n951 NETTRAN_DUMMY_16186 NETTRAN_DUMMY_16187 INV_X32 
XU935 n949 n952 NETTRAN_DUMMY_16188 NETTRAN_DUMMY_16189 INV_X32 
XU936 c0_r2[17] n953 NETTRAN_DUMMY_16190 NETTRAN_DUMMY_16191 CLKBUF_X1 
XU937 n955 n954 NETTRAN_DUMMY_16192 NETTRAN_DUMMY_16193 CLKBUF_X1 
XU938 n953 n955 NETTRAN_DUMMY_16194 NETTRAN_DUMMY_16195 INV_X32 
XU939 n954 n956 NETTRAN_DUMMY_16196 NETTRAN_DUMMY_16197 INV_X32 
XU940 c0_r3[17] n957 NETTRAN_DUMMY_16198 NETTRAN_DUMMY_16199 CLKBUF_X1 
XU941 n959 n958 NETTRAN_DUMMY_16200 NETTRAN_DUMMY_16201 CLKBUF_X1 
XU942 n957 n959 NETTRAN_DUMMY_16202 NETTRAN_DUMMY_16203 INV_X32 
XU943 n958 n960 NETTRAN_DUMMY_16204 NETTRAN_DUMMY_16205 INV_X32 
XU944 c0_r1[16] n961 NETTRAN_DUMMY_16206 NETTRAN_DUMMY_16207 CLKBUF_X1 
XU945 n963 n962 NETTRAN_DUMMY_16208 NETTRAN_DUMMY_16209 CLKBUF_X1 
XU946 n961 n963 NETTRAN_DUMMY_16210 NETTRAN_DUMMY_16211 INV_X32 
XU947 n962 n964 NETTRAN_DUMMY_16212 NETTRAN_DUMMY_16213 INV_X32 
XU948 c0_r2[16] n965 NETTRAN_DUMMY_16214 NETTRAN_DUMMY_16215 CLKBUF_X1 
XU949 n967 n966 NETTRAN_DUMMY_16216 NETTRAN_DUMMY_16217 CLKBUF_X1 
XU950 n965 n967 NETTRAN_DUMMY_16218 NETTRAN_DUMMY_16219 INV_X32 
XU951 n966 n968 NETTRAN_DUMMY_16220 NETTRAN_DUMMY_16221 INV_X32 
XU952 c0_r3[16] n969 NETTRAN_DUMMY_16222 NETTRAN_DUMMY_16223 CLKBUF_X1 
XU953 n971 n970 NETTRAN_DUMMY_16224 NETTRAN_DUMMY_16225 CLKBUF_X1 
XU954 n969 n971 NETTRAN_DUMMY_16226 NETTRAN_DUMMY_16227 INV_X32 
XU955 n970 n972 NETTRAN_DUMMY_16228 NETTRAN_DUMMY_16229 INV_X32 
XU956 c0_r1[15] n973 NETTRAN_DUMMY_16230 NETTRAN_DUMMY_16231 CLKBUF_X1 
XU957 n975 n974 NETTRAN_DUMMY_16232 NETTRAN_DUMMY_16233 CLKBUF_X1 
XU958 n973 n975 NETTRAN_DUMMY_16234 NETTRAN_DUMMY_16235 INV_X32 
XU959 n974 n976 NETTRAN_DUMMY_16236 NETTRAN_DUMMY_16237 INV_X32 
XU960 c0_r2[15] n977 NETTRAN_DUMMY_16238 NETTRAN_DUMMY_16239 CLKBUF_X1 
XU961 n979 n978 NETTRAN_DUMMY_16240 NETTRAN_DUMMY_16241 CLKBUF_X1 
XU962 n977 n979 NETTRAN_DUMMY_16242 NETTRAN_DUMMY_16243 INV_X32 
XU963 n978 n981 NETTRAN_DUMMY_16244 NETTRAN_DUMMY_16245 INV_X32 
XU964 c0_r3[15] n982 NETTRAN_DUMMY_16246 NETTRAN_DUMMY_16247 CLKBUF_X1 
XU965 n984 n983 NETTRAN_DUMMY_16248 NETTRAN_DUMMY_16249 CLKBUF_X1 
XU966 n982 n984 NETTRAN_DUMMY_16250 NETTRAN_DUMMY_16251 INV_X32 
XU967 n983 n985 NETTRAN_DUMMY_16252 NETTRAN_DUMMY_16253 INV_X32 
XU968 c0_r1[14] n986 NETTRAN_DUMMY_16254 NETTRAN_DUMMY_16255 CLKBUF_X1 
XU969 n988 n987 NETTRAN_DUMMY_16256 NETTRAN_DUMMY_16257 CLKBUF_X1 
XU970 n986 n988 NETTRAN_DUMMY_16258 NETTRAN_DUMMY_16259 INV_X32 
XU971 n987 n989 NETTRAN_DUMMY_16260 NETTRAN_DUMMY_16261 INV_X32 
XU972 c0_r2[14] n991 NETTRAN_DUMMY_16262 NETTRAN_DUMMY_16263 CLKBUF_X1 
XU973 n993 n992 NETTRAN_DUMMY_16264 NETTRAN_DUMMY_16265 CLKBUF_X1 
XU974 n991 n993 NETTRAN_DUMMY_16266 NETTRAN_DUMMY_16267 INV_X32 
XU975 n992 n994 NETTRAN_DUMMY_16268 NETTRAN_DUMMY_16269 INV_X32 
XU976 c0_r3[14] n995 NETTRAN_DUMMY_16270 NETTRAN_DUMMY_16271 CLKBUF_X1 
XU977 n997 n996 NETTRAN_DUMMY_16272 NETTRAN_DUMMY_16273 CLKBUF_X1 
XU978 n995 n997 NETTRAN_DUMMY_16274 NETTRAN_DUMMY_16275 INV_X32 
XU979 n996 n998 NETTRAN_DUMMY_16276 NETTRAN_DUMMY_16277 INV_X32 
XU980 c0_r1[13] n999 NETTRAN_DUMMY_16278 NETTRAN_DUMMY_16279 CLKBUF_X1 
XU981 n1002 n1001 NETTRAN_DUMMY_16280 NETTRAN_DUMMY_16281 CLKBUF_X1 
XU982 n999 n1002 NETTRAN_DUMMY_16282 NETTRAN_DUMMY_16283 INV_X32 
XU983 n1001 n1003 NETTRAN_DUMMY_16284 NETTRAN_DUMMY_16285 INV_X32 
XU984 c0_r2[13] n1004 NETTRAN_DUMMY_16286 NETTRAN_DUMMY_16287 CLKBUF_X1 
XU985 n1006 n1005 NETTRAN_DUMMY_16288 NETTRAN_DUMMY_16289 CLKBUF_X1 
XU986 n1004 n1006 NETTRAN_DUMMY_16290 NETTRAN_DUMMY_16291 INV_X32 
XU987 n1005 n1007 NETTRAN_DUMMY_16292 NETTRAN_DUMMY_16293 INV_X32 
XU988 c0_r3[13] n1008 NETTRAN_DUMMY_16294 NETTRAN_DUMMY_16295 CLKBUF_X1 
XU989 n1012 n1009 NETTRAN_DUMMY_16296 NETTRAN_DUMMY_16297 CLKBUF_X1 
XU990 n1008 n1012 NETTRAN_DUMMY_16298 NETTRAN_DUMMY_16299 INV_X32 
XU991 n1009 n1013 NETTRAN_DUMMY_16300 NETTRAN_DUMMY_16301 INV_X32 
XU992 c0_r1[12] n1014 NETTRAN_DUMMY_16302 NETTRAN_DUMMY_16303 CLKBUF_X1 
XU993 n1016 n1015 NETTRAN_DUMMY_16304 NETTRAN_DUMMY_16305 CLKBUF_X1 
XU994 n1014 n1016 NETTRAN_DUMMY_16306 NETTRAN_DUMMY_16307 INV_X32 
XU995 n1015 n1017 NETTRAN_DUMMY_16308 NETTRAN_DUMMY_16309 INV_X32 
XU996 c0_r2[12] n1018 NETTRAN_DUMMY_16310 NETTRAN_DUMMY_16311 CLKBUF_X1 
XU997 n1021 n1019 NETTRAN_DUMMY_16312 NETTRAN_DUMMY_16313 CLKBUF_X1 
XU998 n1018 n1021 NETTRAN_DUMMY_16314 NETTRAN_DUMMY_16315 INV_X32 
XU999 n1019 n1022 NETTRAN_DUMMY_16316 NETTRAN_DUMMY_16317 INV_X32 
XU1000 c0_r3[12] n1023 NETTRAN_DUMMY_16318 NETTRAN_DUMMY_16319 CLKBUF_X1 
XU1001 n1025 n1024 NETTRAN_DUMMY_16320 NETTRAN_DUMMY_16321 CLKBUF_X1 
XU1002 n1023 n1025 NETTRAN_DUMMY_16322 NETTRAN_DUMMY_16323 INV_X32 
XU1003 n1024 n1026 NETTRAN_DUMMY_16324 NETTRAN_DUMMY_16325 INV_X32 
XU1004 c0_r1[11] n1027 NETTRAN_DUMMY_16326 NETTRAN_DUMMY_16327 CLKBUF_X1 
XU1005 n1029 n1028 NETTRAN_DUMMY_16328 NETTRAN_DUMMY_16329 CLKBUF_X1 
XU1006 n1027 n1029 NETTRAN_DUMMY_16330 NETTRAN_DUMMY_16331 INV_X32 
XU1007 n1028 n1031 NETTRAN_DUMMY_16332 NETTRAN_DUMMY_16333 INV_X32 
XU1008 c0_r2[11] n1032 NETTRAN_DUMMY_16334 NETTRAN_DUMMY_16335 CLKBUF_X1 
XU1009 n1034 n1033 NETTRAN_DUMMY_16336 NETTRAN_DUMMY_16337 CLKBUF_X1 
XU1010 n1032 n1034 NETTRAN_DUMMY_16338 NETTRAN_DUMMY_16339 INV_X32 
XU1011 n1033 n1035 NETTRAN_DUMMY_16340 NETTRAN_DUMMY_16341 INV_X32 
XU1012 c0_r3[11] n1036 NETTRAN_DUMMY_16342 NETTRAN_DUMMY_16343 CLKBUF_X1 
XU1013 n1038 n1037 NETTRAN_DUMMY_16344 NETTRAN_DUMMY_16345 CLKBUF_X1 
XU1014 n1036 n1038 NETTRAN_DUMMY_16346 NETTRAN_DUMMY_16347 INV_X32 
XU1015 n1037 n1039 NETTRAN_DUMMY_16348 NETTRAN_DUMMY_16349 INV_X32 
XU1016 c0_r1[10] n1041 NETTRAN_DUMMY_16350 NETTRAN_DUMMY_16351 CLKBUF_X1 
XU1017 n1043 n1042 NETTRAN_DUMMY_16352 NETTRAN_DUMMY_16353 CLKBUF_X1 
XU1018 n1041 n1043 NETTRAN_DUMMY_16354 NETTRAN_DUMMY_16355 INV_X32 
XU1019 n1042 n1044 NETTRAN_DUMMY_16356 NETTRAN_DUMMY_16357 INV_X32 
XU1020 c0_r2[10] n1045 NETTRAN_DUMMY_16358 NETTRAN_DUMMY_16359 CLKBUF_X1 
XU1021 n1047 n1046 NETTRAN_DUMMY_16360 NETTRAN_DUMMY_16361 CLKBUF_X1 
XU1022 n1045 n1047 NETTRAN_DUMMY_16362 NETTRAN_DUMMY_16363 INV_X32 
XU1023 n1046 n1048 NETTRAN_DUMMY_16364 NETTRAN_DUMMY_16365 INV_X32 
XU1024 n1053 n1049 NETTRAN_DUMMY_16366 NETTRAN_DUMMY_16367 BUF_X1 
XU1025 n1052 n1051 NETTRAN_DUMMY_16368 NETTRAN_DUMMY_16369 CLKBUF_X1 
XU1026 c0_r3[10] n1052 NETTRAN_DUMMY_16370 NETTRAN_DUMMY_16371 INV_X32 
XU1027 n1051 n1053 NETTRAN_DUMMY_16372 NETTRAN_DUMMY_16373 INV_X32 
XU1028 c0_r1[9] n1054 NETTRAN_DUMMY_16374 NETTRAN_DUMMY_16375 CLKBUF_X1 
XU1029 n1900 n1055 NETTRAN_DUMMY_16376 NETTRAN_DUMMY_16377 CLKBUF_X1 
XU1030 n1054 n1056 NETTRAN_DUMMY_16378 NETTRAN_DUMMY_16379 INV_X32 
XU1031 n1055 n1057 NETTRAN_DUMMY_16380 NETTRAN_DUMMY_16381 INV_X32 
XU1032 c0_r2[9] n1058 NETTRAN_DUMMY_16382 NETTRAN_DUMMY_16383 CLKBUF_X1 
XU1033 n1061 n1059 NETTRAN_DUMMY_16384 NETTRAN_DUMMY_16385 CLKBUF_X1 
XU1034 n1058 n1061 NETTRAN_DUMMY_16386 NETTRAN_DUMMY_16387 INV_X32 
XU1035 n1059 n1062 NETTRAN_DUMMY_16388 NETTRAN_DUMMY_16389 INV_X32 
XU1036 c0_r3[9] n1063 NETTRAN_DUMMY_16390 NETTRAN_DUMMY_16391 CLKBUF_X1 
XU1037 n1065 n1064 NETTRAN_DUMMY_16392 NETTRAN_DUMMY_16393 CLKBUF_X1 
XU1038 n1063 n1065 NETTRAN_DUMMY_16394 NETTRAN_DUMMY_16395 INV_X32 
XU1039 n1064 n1066 NETTRAN_DUMMY_16396 NETTRAN_DUMMY_16397 INV_X32 
XU1040 c0_r1[8] n1067 NETTRAN_DUMMY_16398 NETTRAN_DUMMY_16399 CLKBUF_X1 
XU1041 n1069 n1068 NETTRAN_DUMMY_16400 NETTRAN_DUMMY_16401 CLKBUF_X1 
XU1042 n1067 n1069 NETTRAN_DUMMY_16402 NETTRAN_DUMMY_16403 INV_X32 
XU1043 n1068 n1071 NETTRAN_DUMMY_16404 NETTRAN_DUMMY_16405 INV_X32 
XU1044 N11000 n1072 NETTRAN_DUMMY_16406 NETTRAN_DUMMY_16407 INV_X1 
XU1045 n1072 n1073 NETTRAN_DUMMY_16408 NETTRAN_DUMMY_16409 INV_X32 
XU1046 n1077 n1074 NETTRAN_DUMMY_16410 NETTRAN_DUMMY_16411 INV_X1 
XU1047 n1074 n1075 NETTRAN_DUMMY_16412 NETTRAN_DUMMY_16413 INV_X32 
XU1048 N10 n1076 NETTRAN_DUMMY_16414 NETTRAN_DUMMY_16415 INV_X1 
XU1049 n1076 n1077 NETTRAN_DUMMY_16416 NETTRAN_DUMMY_16417 INV_X32 
XU1050 N900 n1078 NETTRAN_DUMMY_16418 NETTRAN_DUMMY_16419 INV_X1 
XU1051 n1078 n1079 NETTRAN_DUMMY_16420 NETTRAN_DUMMY_16421 INV_X32 
XU1052 N8 n1081 NETTRAN_DUMMY_16422 NETTRAN_DUMMY_16423 BUF_X1 
XU1053 N700 n1082 NETTRAN_DUMMY_16424 NETTRAN_DUMMY_16425 CLKBUF_X1 
XU1054 N74 n1083 NETTRAN_DUMMY_16426 NETTRAN_DUMMY_16427 CLKBUF_X1 
XU1055 n1117 n1084 NETTRAN_DUMMY_16428 NETTRAN_DUMMY_16429 BUF_X1 
XU1056 N7010 n1085 NETTRAN_DUMMY_16430 NETTRAN_DUMMY_16431 BUF_X1 
XU1057 n7210 n1086 NETTRAN_DUMMY_16432 NETTRAN_DUMMY_16433 BUF_X1 
XU1058 num_lzd_r[3] n1087 NETTRAN_DUMMY_16434 NETTRAN_DUMMY_16435 INV_X1 
XU1059 n1087 n1088 NETTRAN_DUMMY_16436 NETTRAN_DUMMY_16437 INV_X32 
XU1060 n1010 n1089 NETTRAN_DUMMY_16438 NETTRAN_DUMMY_16439 INV_X1 
XU1061 n1089 n1091 NETTRAN_DUMMY_16440 NETTRAN_DUMMY_16441 INV_X32 
XU1062 n205 n10921 NETTRAN_DUMMY_16442 NETTRAN_DUMMY_16443 CLKBUF_X1 
XU1063 n810 n1093 NETTRAN_DUMMY_16444 NETTRAN_DUMMY_16445 CLKBUF_X1 
XU1064 n1110 n1094 NETTRAN_DUMMY_16446 NETTRAN_DUMMY_16447 INV_X1 
XU1065 n1094 n1095 NETTRAN_DUMMY_16448 NETTRAN_DUMMY_16449 INV_X16 
XU1066 n143 n1096 NETTRAN_DUMMY_16450 NETTRAN_DUMMY_16451 CLKBUF_X1 
XU1067 num_lzd_r[5] n1097 NETTRAN_DUMMY_16452 NETTRAN_DUMMY_16453 INV_X1 
XU1068 n1097 n1098 NETTRAN_DUMMY_16454 NETTRAN_DUMMY_16455 INV_X32 
XU1069 num_lzd_r[4] n1099 NETTRAN_DUMMY_16456 NETTRAN_DUMMY_16457 INV_X32 
XU1070 n1099 n1101 NETTRAN_DUMMY_16458 NETTRAN_DUMMY_16459 INV_X1 
XU1071 N65 n1102 NETTRAN_DUMMY_16460 NETTRAN_DUMMY_16461 INV_X1 
XU1072 n46 n1104 NETTRAN_DUMMY_16462 NETTRAN_DUMMY_16463 INV_X1 
XU1073 n1104 n1105 NETTRAN_DUMMY_16464 NETTRAN_DUMMY_16465 INV_X32 
XU1074 n1105 n1106 NETTRAN_DUMMY_16466 NETTRAN_DUMMY_16467 INV_X1 
XU1075 n1106 n1107 NETTRAN_DUMMY_16468 NETTRAN_DUMMY_16469 INV_X32 
XU1076 N64 n1108 NETTRAN_DUMMY_16470 NETTRAN_DUMMY_16471 INV_X1 
XU1077 n48 n1112 NETTRAN_DUMMY_16472 NETTRAN_DUMMY_16473 INV_X1 
XU1078 n1112 n1113 NETTRAN_DUMMY_16474 NETTRAN_DUMMY_16475 INV_X32 
XU1079 n1113 n1114 NETTRAN_DUMMY_16476 NETTRAN_DUMMY_16477 INV_X1 
XU1080 n1114 n1115 NETTRAN_DUMMY_16478 NETTRAN_DUMMY_16479 INV_X32 
XU1081 n50 n1116 NETTRAN_DUMMY_16480 NETTRAN_DUMMY_16481 INV_X32 
XU1082 n1122 n1118 NETTRAN_DUMMY_16482 NETTRAN_DUMMY_16483 INV_X1 
XU1083 n1118 n1119 NETTRAN_DUMMY_16484 NETTRAN_DUMMY_16485 INV_X32 
XU1084 n49 n1121 NETTRAN_DUMMY_16486 NETTRAN_DUMMY_16487 INV_X1 
XU1085 n1121 n1122 NETTRAN_DUMMY_16488 NETTRAN_DUMMY_16489 INV_X32 
XU1086 n1126 n1123 NETTRAN_DUMMY_16490 NETTRAN_DUMMY_16491 CLKBUF_X1 
XU1087 n910 n1124 NETTRAN_DUMMY_16492 NETTRAN_DUMMY_16493 INV_X1 
XU1088 n1124 n1125 NETTRAN_DUMMY_16494 NETTRAN_DUMMY_16495 INV_X32 
XU1089 n1093 n1126 NETTRAN_DUMMY_16496 NETTRAN_DUMMY_16497 INV_X32 
XU1090 N611 n1128 NETTRAN_DUMMY_16498 NETTRAN_DUMMY_16499 INV_X1 
XU1091 n1128 n1129 NETTRAN_DUMMY_16500 NETTRAN_DUMMY_16501 INV_X16 
XU1092 n53 n1130 NETTRAN_DUMMY_16502 NETTRAN_DUMMY_16503 INV_X1 
XU1093 n1130 n1131 NETTRAN_DUMMY_16504 NETTRAN_DUMMY_16505 INV_X32 
XU1094 n1131 n1132 NETTRAN_DUMMY_16506 NETTRAN_DUMMY_16507 INV_X1 
XU1095 n1132 n1133 NETTRAN_DUMMY_16508 NETTRAN_DUMMY_16509 INV_X32 
XU1096 n1137 n1134 NETTRAN_DUMMY_16510 NETTRAN_DUMMY_16511 BUF_X1 
XU1097 n1136 n1135 NETTRAN_DUMMY_16512 NETTRAN_DUMMY_16513 CLKBUF_X1 
XU1098 N600 n1136 NETTRAN_DUMMY_16514 NETTRAN_DUMMY_16515 INV_X32 
XU1099 n1135 n1137 NETTRAN_DUMMY_16516 NETTRAN_DUMMY_16517 INV_X32 
XU1100 N76 n1138 NETTRAN_DUMMY_16518 NETTRAN_DUMMY_16519 CLKBUF_X1 
XU1101 n1140 n1139 NETTRAN_DUMMY_16520 NETTRAN_DUMMY_16521 CLKBUF_X1 
XU1102 n1138 n1140 NETTRAN_DUMMY_16522 NETTRAN_DUMMY_16523 INV_X32 
XU1103 n1139 n1141 NETTRAN_DUMMY_16524 NETTRAN_DUMMY_16525 INV_X32 
XU1104 n1145 n1142 NETTRAN_DUMMY_16526 NETTRAN_DUMMY_16527 BUF_X1 
XU1105 n1144 n1143 NETTRAN_DUMMY_16528 NETTRAN_DUMMY_16529 CLKBUF_X1 
XU1106 N75 n1144 NETTRAN_DUMMY_16530 NETTRAN_DUMMY_16531 INV_X32 
XU1107 n1143 n1145 NETTRAN_DUMMY_16532 NETTRAN_DUMMY_16533 INV_X32 
XU1108 N91 n1146 NETTRAN_DUMMY_16534 NETTRAN_DUMMY_16535 CLKBUF_X1 
XU1109 n1148 n1147 NETTRAN_DUMMY_16536 NETTRAN_DUMMY_16537 CLKBUF_X1 
XU1110 n1146 n1148 NETTRAN_DUMMY_16538 NETTRAN_DUMMY_16539 INV_X32 
XU1111 n1147 n1149 NETTRAN_DUMMY_16540 NETTRAN_DUMMY_16541 INV_X32 
XU1112 N9010 n1150 NETTRAN_DUMMY_16542 NETTRAN_DUMMY_16543 CLKBUF_X1 
XU1113 n1152 n1151 NETTRAN_DUMMY_16544 NETTRAN_DUMMY_16545 CLKBUF_X1 
XU1114 n1150 n1152 NETTRAN_DUMMY_16546 NETTRAN_DUMMY_16547 INV_X32 
XU1115 n1151 n1153 NETTRAN_DUMMY_16548 NETTRAN_DUMMY_16549 INV_X32 
XU1116 N89 n1154 NETTRAN_DUMMY_16550 NETTRAN_DUMMY_16551 CLKBUF_X1 
XU1117 n1156 n1155 NETTRAN_DUMMY_16552 NETTRAN_DUMMY_16553 CLKBUF_X1 
XU1118 n1154 n1156 NETTRAN_DUMMY_16554 NETTRAN_DUMMY_16555 INV_X32 
XU1119 n1155 n1157 NETTRAN_DUMMY_16556 NETTRAN_DUMMY_16557 INV_X32 
XU1120 N88 n1158 NETTRAN_DUMMY_16558 NETTRAN_DUMMY_16559 INV_X1 
XU1121 n1930 n1159 NETTRAN_DUMMY_16560 NETTRAN_DUMMY_16561 INV_X32 
XU1122 N87 n1160 NETTRAN_DUMMY_16562 NETTRAN_DUMMY_16563 CLKBUF_X1 
XU1123 n1162 n1161 NETTRAN_DUMMY_16564 NETTRAN_DUMMY_16565 CLKBUF_X1 
XU1124 n1160 n1162 NETTRAN_DUMMY_16566 NETTRAN_DUMMY_16567 INV_X32 
XU1125 n1161 n1163 NETTRAN_DUMMY_16568 NETTRAN_DUMMY_16569 INV_X32 
XU1126 n1165 n1164 NETTRAN_DUMMY_16570 NETTRAN_DUMMY_16571 CLKBUF_X1 
XU1127 N86 n1165 NETTRAN_DUMMY_16572 NETTRAN_DUMMY_16573 INV_X32 
XU1128 n1164 n1166 NETTRAN_DUMMY_16574 NETTRAN_DUMMY_16575 INV_X32 
XU1129 n1170 n1167 NETTRAN_DUMMY_16576 NETTRAN_DUMMY_16577 CLKBUF_X1 
XU1130 n1169 n1168 NETTRAN_DUMMY_16578 NETTRAN_DUMMY_16579 CLKBUF_X1 
XU1131 N85 n1169 NETTRAN_DUMMY_16580 NETTRAN_DUMMY_16581 INV_X32 
XU1132 n1168 n1170 NETTRAN_DUMMY_16582 NETTRAN_DUMMY_16583 INV_X32 
XU1133 N84 n1171 NETTRAN_DUMMY_16584 NETTRAN_DUMMY_16585 CLKBUF_X1 
XU1134 n1173 n1172 NETTRAN_DUMMY_16586 NETTRAN_DUMMY_16587 CLKBUF_X1 
XU1135 n1171 n1173 NETTRAN_DUMMY_16588 NETTRAN_DUMMY_16589 INV_X32 
XU1136 n1172 n1174 NETTRAN_DUMMY_16590 NETTRAN_DUMMY_16591 INV_X32 
XU1137 N83 n1175 NETTRAN_DUMMY_16592 NETTRAN_DUMMY_16593 CLKBUF_X1 
XU1138 n1177 n1176 NETTRAN_DUMMY_16594 NETTRAN_DUMMY_16595 CLKBUF_X1 
XU1139 n1175 n1177 NETTRAN_DUMMY_16596 NETTRAN_DUMMY_16597 INV_X32 
XU1140 n1176 n1178 NETTRAN_DUMMY_16598 NETTRAN_DUMMY_16599 INV_X32 
XU1141 N82 n1179 NETTRAN_DUMMY_16600 NETTRAN_DUMMY_16601 CLKBUF_X1 
XU1142 n1181 n1180 NETTRAN_DUMMY_16602 NETTRAN_DUMMY_16603 CLKBUF_X1 
XU1143 n1179 n1181 NETTRAN_DUMMY_16604 NETTRAN_DUMMY_16605 INV_X32 
XU1144 n1180 n1182 NETTRAN_DUMMY_16606 NETTRAN_DUMMY_16607 INV_X32 
XU1145 N81 n1183 NETTRAN_DUMMY_16608 NETTRAN_DUMMY_16609 CLKBUF_X1 
XU1146 n1185 n1184 NETTRAN_DUMMY_16610 NETTRAN_DUMMY_16611 CLKBUF_X1 
XU1147 n1183 n1185 NETTRAN_DUMMY_16612 NETTRAN_DUMMY_16613 INV_X32 
XU1148 n1184 n1186 NETTRAN_DUMMY_16614 NETTRAN_DUMMY_16615 INV_X32 
XU1149 N79 n1187 NETTRAN_DUMMY_16616 NETTRAN_DUMMY_16617 CLKBUF_X1 
XU1150 n1189 n1188 NETTRAN_DUMMY_16618 NETTRAN_DUMMY_16619 CLKBUF_X1 
XU1151 n1187 n1189 NETTRAN_DUMMY_16620 NETTRAN_DUMMY_16621 INV_X32 
XU1152 n1188 n1190 NETTRAN_DUMMY_16622 NETTRAN_DUMMY_16623 INV_X32 
XU1153 n1194 n1191 NETTRAN_DUMMY_16624 NETTRAN_DUMMY_16625 BUF_X1 
XU1154 n1193 n1192 NETTRAN_DUMMY_16626 NETTRAN_DUMMY_16627 CLKBUF_X1 
XU1155 N78 n1193 NETTRAN_DUMMY_16628 NETTRAN_DUMMY_16629 INV_X32 
XU1156 n1192 n1194 NETTRAN_DUMMY_16630 NETTRAN_DUMMY_16631 INV_X32 
XU1157 n1198 n1195 NETTRAN_DUMMY_16632 NETTRAN_DUMMY_16633 BUF_X1 
XU1158 n1197 n1196 NETTRAN_DUMMY_16634 NETTRAN_DUMMY_16635 CLKBUF_X1 
XU1159 N77 n1197 NETTRAN_DUMMY_16636 NETTRAN_DUMMY_16637 INV_X32 
XU1160 n1196 n1198 NETTRAN_DUMMY_16638 NETTRAN_DUMMY_16639 INV_X32 
XU1161 n1201 n1199 NETTRAN_DUMMY_16640 NETTRAN_DUMMY_16641 INV_X32 
XU1162 n1199 n1200 NETTRAN_DUMMY_16642 NETTRAN_DUMMY_16643 INV_X1 
XU1163 n1204 n1201 NETTRAN_DUMMY_16644 NETTRAN_DUMMY_16645 INV_X1 
XU1164 n1200 n1202 NETTRAN_DUMMY_16646 NETTRAN_DUMMY_16647 INV_X32 
XU1165 N92 n1203 NETTRAN_DUMMY_16648 NETTRAN_DUMMY_16649 INV_X1 
XU1166 n1203 n1204 NETTRAN_DUMMY_16650 NETTRAN_DUMMY_16651 INV_X32 
XU1167 x_r1[14] n1205 NETTRAN_DUMMY_16652 NETTRAN_DUMMY_16653 CLKBUF_X1 
XU1168 n1207 n1206 NETTRAN_DUMMY_16654 NETTRAN_DUMMY_16655 CLKBUF_X1 
XU1169 n1205 n1207 NETTRAN_DUMMY_16656 NETTRAN_DUMMY_16657 INV_X32 
XU1170 n1206 n1208 NETTRAN_DUMMY_16658 NETTRAN_DUMMY_16659 INV_X32 
XU1171 x_r2[14] n1209 NETTRAN_DUMMY_16660 NETTRAN_DUMMY_16661 CLKBUF_X1 
XU1172 n1211 n1210 NETTRAN_DUMMY_16662 NETTRAN_DUMMY_16663 CLKBUF_X1 
XU1173 n1209 n1211 NETTRAN_DUMMY_16664 NETTRAN_DUMMY_16665 INV_X32 
XU1174 n1210 n1212 NETTRAN_DUMMY_16666 NETTRAN_DUMMY_16667 INV_X32 
XU1175 n1215 n1213 NETTRAN_DUMMY_16668 NETTRAN_DUMMY_16669 INV_X32 
XU1176 n1213 n1214 NETTRAN_DUMMY_16670 NETTRAN_DUMMY_16671 INV_X1 
XU1177 n1218 n1215 NETTRAN_DUMMY_16672 NETTRAN_DUMMY_16673 INV_X1 
XU1178 n1214 n1216 NETTRAN_DUMMY_16674 NETTRAN_DUMMY_16675 INV_X32 
XU1179 N93 n1217 NETTRAN_DUMMY_16676 NETTRAN_DUMMY_16677 INV_X1 
XU1180 n1217 n1218 NETTRAN_DUMMY_16678 NETTRAN_DUMMY_16679 INV_X32 
XU1181 x_r1[13] n1219 NETTRAN_DUMMY_16680 NETTRAN_DUMMY_16681 CLKBUF_X1 
XU1182 n1221 n1220 NETTRAN_DUMMY_16682 NETTRAN_DUMMY_16683 CLKBUF_X1 
XU1183 n1219 n1221 NETTRAN_DUMMY_16684 NETTRAN_DUMMY_16685 INV_X32 
XU1184 n1220 n1222 NETTRAN_DUMMY_16686 NETTRAN_DUMMY_16687 INV_X32 
XU1185 x_r2[13] n1223 NETTRAN_DUMMY_16688 NETTRAN_DUMMY_16689 CLKBUF_X1 
XU1186 n1225 n1224 NETTRAN_DUMMY_16690 NETTRAN_DUMMY_16691 CLKBUF_X1 
XU1187 n1223 n1225 NETTRAN_DUMMY_16692 NETTRAN_DUMMY_16693 INV_X32 
XU1188 n1224 n1226 NETTRAN_DUMMY_16694 NETTRAN_DUMMY_16695 INV_X32 
XU1189 n1228 n1227 NETTRAN_DUMMY_16696 NETTRAN_DUMMY_16697 CLKBUF_X1 
XU1190 n1231 n1228 NETTRAN_DUMMY_16698 NETTRAN_DUMMY_16699 INV_X1 
XU1191 n1227 n1229 NETTRAN_DUMMY_16700 NETTRAN_DUMMY_16701 INV_X32 
XU1192 N94 n1230 NETTRAN_DUMMY_16702 NETTRAN_DUMMY_16703 INV_X1 
XU1193 n1230 n1231 NETTRAN_DUMMY_16704 NETTRAN_DUMMY_16705 INV_X32 
XU1194 x_r1[12] n1232 NETTRAN_DUMMY_16706 NETTRAN_DUMMY_16707 CLKBUF_X1 
XU1195 n1234 n1233 NETTRAN_DUMMY_16708 NETTRAN_DUMMY_16709 CLKBUF_X1 
XU1196 n1232 n1234 NETTRAN_DUMMY_16710 NETTRAN_DUMMY_16711 INV_X32 
XU1197 n1233 n1235 NETTRAN_DUMMY_16712 NETTRAN_DUMMY_16713 INV_X32 
XU1198 x_r2[12] n1236 NETTRAN_DUMMY_16714 NETTRAN_DUMMY_16715 CLKBUF_X1 
XU1199 n1238 n1237 NETTRAN_DUMMY_16716 NETTRAN_DUMMY_16717 CLKBUF_X1 
XU1200 n1236 n1238 NETTRAN_DUMMY_16718 NETTRAN_DUMMY_16719 INV_X32 
XU1201 n1237 n1239 NETTRAN_DUMMY_16720 NETTRAN_DUMMY_16721 INV_X32 
XU1202 n1242 n1240 NETTRAN_DUMMY_16722 NETTRAN_DUMMY_16723 INV_X32 
XU1203 n1240 n1241 NETTRAN_DUMMY_16724 NETTRAN_DUMMY_16725 INV_X1 
XU1204 N95 n1242 NETTRAN_DUMMY_16726 NETTRAN_DUMMY_16727 INV_X1 
XU1205 n1241 n1243 NETTRAN_DUMMY_16728 NETTRAN_DUMMY_16729 INV_X32 
XU1206 n1243 n1244 NETTRAN_DUMMY_16730 NETTRAN_DUMMY_16731 INV_X1 
XU1207 n1244 n1245 NETTRAN_DUMMY_16732 NETTRAN_DUMMY_16733 INV_X32 
XU1208 x_r1[11] n1246 NETTRAN_DUMMY_16734 NETTRAN_DUMMY_16735 CLKBUF_X1 
XU1209 n1248 n1247 NETTRAN_DUMMY_16736 NETTRAN_DUMMY_16737 CLKBUF_X1 
XU1210 n1246 n1248 NETTRAN_DUMMY_16738 NETTRAN_DUMMY_16739 INV_X32 
XU1211 n1247 n1249 NETTRAN_DUMMY_16740 NETTRAN_DUMMY_16741 INV_X32 
XU1212 x_r2[11] n1250 NETTRAN_DUMMY_16742 NETTRAN_DUMMY_16743 CLKBUF_X1 
XU1213 n1252 n1251 NETTRAN_DUMMY_16744 NETTRAN_DUMMY_16745 CLKBUF_X1 
XU1214 n1250 n1252 NETTRAN_DUMMY_16746 NETTRAN_DUMMY_16747 INV_X32 
XU1215 n1251 n1253 NETTRAN_DUMMY_16748 NETTRAN_DUMMY_16749 INV_X32 
XU1216 n1255 n1254 NETTRAN_DUMMY_16750 NETTRAN_DUMMY_16751 CLKBUF_X1 
XU1217 N96 n1255 NETTRAN_DUMMY_16752 NETTRAN_DUMMY_16753 INV_X1 
XU1218 n1254 n1256 NETTRAN_DUMMY_16754 NETTRAN_DUMMY_16755 INV_X32 
XU1219 n1256 n1257 NETTRAN_DUMMY_16756 NETTRAN_DUMMY_16757 INV_X1 
XU1220 n1257 n1258 NETTRAN_DUMMY_16758 NETTRAN_DUMMY_16759 INV_X32 
XU1221 x_r1[10] n1259 NETTRAN_DUMMY_16760 NETTRAN_DUMMY_16761 CLKBUF_X1 
XU1222 n1261 n1260 NETTRAN_DUMMY_16762 NETTRAN_DUMMY_16763 CLKBUF_X1 
XU1223 n1259 n1261 NETTRAN_DUMMY_16764 NETTRAN_DUMMY_16765 INV_X32 
XU1224 n1260 n1262 NETTRAN_DUMMY_16766 NETTRAN_DUMMY_16767 INV_X32 
XU1225 x_r2[10] n1263 NETTRAN_DUMMY_16768 NETTRAN_DUMMY_16769 CLKBUF_X1 
XU1226 n1265 n1264 NETTRAN_DUMMY_16770 NETTRAN_DUMMY_16771 CLKBUF_X1 
XU1227 n1263 n1265 NETTRAN_DUMMY_16772 NETTRAN_DUMMY_16773 INV_X32 
XU1228 n1264 n1266 NETTRAN_DUMMY_16774 NETTRAN_DUMMY_16775 INV_X32 
XU1229 n1270 n1267 NETTRAN_DUMMY_16776 NETTRAN_DUMMY_16777 INV_X1 
XU1231 n1272 n1269 NETTRAN_DUMMY_16778 NETTRAN_DUMMY_16779 INV_X1 
XU1232 n1269 n1270 NETTRAN_DUMMY_16780 NETTRAN_DUMMY_16781 INV_X32 
XU1233 N97 n1271 NETTRAN_DUMMY_16782 NETTRAN_DUMMY_16783 INV_X1 
XU1234 n1271 n1272 NETTRAN_DUMMY_16784 NETTRAN_DUMMY_16785 INV_X32 
XU1235 x_r1[9] n1273 NETTRAN_DUMMY_16786 NETTRAN_DUMMY_16787 CLKBUF_X1 
XU1236 n1275 n1274 NETTRAN_DUMMY_16788 NETTRAN_DUMMY_16789 CLKBUF_X1 
XU1237 n1273 n1275 NETTRAN_DUMMY_16790 NETTRAN_DUMMY_16791 INV_X32 
XU1238 n1274 n1276 NETTRAN_DUMMY_16792 NETTRAN_DUMMY_16793 INV_X32 
XU1239 x_r2[9] n1277 NETTRAN_DUMMY_16794 NETTRAN_DUMMY_16795 CLKBUF_X1 
XU1240 n1279 n1278 NETTRAN_DUMMY_16796 NETTRAN_DUMMY_16797 CLKBUF_X1 
XU1241 n1277 n1279 NETTRAN_DUMMY_16798 NETTRAN_DUMMY_16799 INV_X32 
XU1242 n1278 n1280 NETTRAN_DUMMY_16800 NETTRAN_DUMMY_16801 INV_X32 
XU1243 n1284 n1281 NETTRAN_DUMMY_16802 NETTRAN_DUMMY_16803 CLKBUF_X1 
XU1244 N98 n1282 NETTRAN_DUMMY_16804 NETTRAN_DUMMY_16805 INV_X1 
XU1245 n1282 n1283 NETTRAN_DUMMY_16806 NETTRAN_DUMMY_16807 INV_X32 
XU1246 n1283 n1284 NETTRAN_DUMMY_16808 NETTRAN_DUMMY_16809 INV_X1 
XU1247 n1281 n1285 NETTRAN_DUMMY_16810 NETTRAN_DUMMY_16811 INV_X32 
XU1248 x_r1[8] n1286 NETTRAN_DUMMY_16812 NETTRAN_DUMMY_16813 CLKBUF_X1 
XU1249 n1288 n1287 NETTRAN_DUMMY_16814 NETTRAN_DUMMY_16815 CLKBUF_X1 
XU1250 n1286 n1288 NETTRAN_DUMMY_16816 NETTRAN_DUMMY_16817 INV_X32 
XU1251 n1287 n1289 NETTRAN_DUMMY_16818 NETTRAN_DUMMY_16819 INV_X32 
XU1252 x_r2[8] n1290 NETTRAN_DUMMY_16820 NETTRAN_DUMMY_16821 CLKBUF_X1 
XU1253 n1292 n1291 NETTRAN_DUMMY_16822 NETTRAN_DUMMY_16823 CLKBUF_X1 
XU1254 n1290 n1292 NETTRAN_DUMMY_16824 NETTRAN_DUMMY_16825 INV_X32 
XU1255 n1291 n1293 NETTRAN_DUMMY_16826 NETTRAN_DUMMY_16827 INV_X32 
XU1256 n1298 n1294 NETTRAN_DUMMY_16828 NETTRAN_DUMMY_16829 INV_X32 
XU1257 n1294 n1295 NETTRAN_DUMMY_16830 NETTRAN_DUMMY_16831 INV_X1 
XU1258 N99 n1296 NETTRAN_DUMMY_16832 NETTRAN_DUMMY_16833 INV_X1 
XU1259 n1296 n1297 NETTRAN_DUMMY_16834 NETTRAN_DUMMY_16835 INV_X32 
XU1260 n1297 n1298 NETTRAN_DUMMY_16836 NETTRAN_DUMMY_16837 INV_X1 
XU1261 n1295 n1299 NETTRAN_DUMMY_16838 NETTRAN_DUMMY_16839 INV_X32 
XU1262 x_r1[7] n1300 NETTRAN_DUMMY_16840 NETTRAN_DUMMY_16841 CLKBUF_X1 
XU1263 n1302 n1301 NETTRAN_DUMMY_16842 NETTRAN_DUMMY_16843 CLKBUF_X1 
XU1264 n1300 n1302 NETTRAN_DUMMY_16844 NETTRAN_DUMMY_16845 INV_X32 
XU1265 n1301 n1303 NETTRAN_DUMMY_16846 NETTRAN_DUMMY_16847 INV_X32 
XU1230 n1267 n1268 NETTRAN_DUMMY_16848 NETTRAN_DUMMY_16849 INV_X16 
XU1266 n446 n1304 NETTRAN_DUMMY_16850 NETTRAN_DUMMY_16851 BUF_X1 
XU1267 N127 n1305 NETTRAN_DUMMY_16852 NETTRAN_DUMMY_16853 BUF_X1 
XU1268 n1268 n1306 NETTRAN_DUMMY_16854 NETTRAN_DUMMY_16855 BUF_X1 
XU1269 n1306 n1307 NETTRAN_DUMMY_16856 NETTRAN_DUMMY_16857 BUF_X1 
XU1294 n135 n1332 NETTRAN_DUMMY_16858 NETTRAN_DUMMY_16859 BUF_X1 
XU1295 n425 n1333 NETTRAN_DUMMY_16860 NETTRAN_DUMMY_16861 BUF_X1 
XU1296 n1285 n1334 NETTRAN_DUMMY_16862 NETTRAN_DUMMY_16863 BUF_X1 
XU1270 N121 n1335 NETTRAN_DUMMY_16864 NETTRAN_DUMMY_16865 BUF_X1 
XU1271 n1335 n1336 NETTRAN_DUMMY_16866 NETTRAN_DUMMY_16867 BUF_X1 
Xu_gng_lzd num_lzd[5] num_lzd[4] num_lzd[3] num_lzd[2] num_lzd[1] num_lzd[0] data_in[63] 
+ data_in[62] data_in[61] data_in[60] data_in[59] data_in[58] data_in[57] data_in[56] 
+ data_in[55] data_in[54] data_in[53] data_in[52] data_in[51] data_in[50] data_in[49] 
+ data_in[48] data_in[47] data_in[46] data_in[45] data_in[44] data_in[43] data_in[42] 
+ data_in[41] data_in[40] data_in[39] data_in[38] data_in[37] data_in[36] data_in[35] 
+ data_in[34] data_in[33] data_in[32] data_in[31] data_in[30] data_in[29] data_in[28] 
+ data_in[27] data_in[26] data_in[25] data_in[24] data_in[23] data_in[22] data_in[21] 
+ data_in[20] data_in[19] data_in[18] data_in[17] data_in[16] data_in[15] data_in[14] 
+ data_in[13] data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] data_in[7] 
+ data_in[6] data_in[5] data_in[4] data_in[3] gng_lzd 
Xu_gng_coef c2[16] c2[15] c2[14] c2[13] c2[12] c2[11] c2[10] c2[9] c2[8] c2[7] c2[6] 
+ c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] n6310 c1[17] c1[16] c1[15] c1[14] c1[13] c1[12] 
+ c1[11] c1[10] c1[9] c1[8] c1[7] c1[6] c1[5] c1[4] c1[3] c1[2] c1[1] c1[0] c0[17] 
+ c0[16] c0[15] c0[14] c0[13] c0[12] c0[11] c0[10] c0[9] c0[8] c0[7] c0[6] c0[5] 
+ c0[4] c0[3] c0[2] c0[1] c0[0] n6810 n10921 n7011 n1096 n7210 n7310 n202 n207 n132 
+ n133 n143 n142 n205 n1332 n63_G2B1I8 n63_G2B1I2 gng_coef 
Xu_gng_smul_16_18_sadd_37 sum1[37] sum1[36] sum1[35] sum1[34] sum1[33] sum1[32] 
+ sum1[31] sum1[30] sum1[29] sum1[28] sum1[27] sum1[26] sum1[25] sum1[24] sum1[23] 
+ sum1[22] sum1[21] sum1[20] SYNOPSYS_UNCONNECTED_26 SYNOPSYS_UNCONNECTED_25 SYNOPSYS_UNCONNECTED_24 
+ SYNOPSYS_UNCONNECTED_34 SYNOPSYS_UNCONNECTED_33 SYNOPSYS_UNCONNECTED_32 SYNOPSYS_UNCONNECTED_31 
+ SYNOPSYS_UNCONNECTED_30 SYNOPSYS_UNCONNECTED_29 SYNOPSYS_UNCONNECTED_28 SYNOPSYS_UNCONNECTED_27 
+ SYNOPSYS_UNCONNECTED_42 SYNOPSYS_UNCONNECTED_41 SYNOPSYS_UNCONNECTED_40 SYNOPSYS_UNCONNECTED_39 
+ SYNOPSYS_UNCONNECTED_38 SYNOPSYS_UNCONNECTED_37 SYNOPSYS_UNCONNECTED_36 SYNOPSYS_UNCONNECTED_35 
+ SYNOPSYS_UNCONNECTED_43 n10920 n214 n218 n222 n226 n230 n234 n145 n242 n246 n250 
+ n1470 n258 n262 n266 n270 n148 n278 n282 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS c2[16] c2[15] c2[14] c2[13] c2[12] c2[11] 
+ c2[10] c2[9] c2[8] c2[7] c2[6] c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] VSS n1208 n1222 
+ n1235 n1249 n1262 n1276 n209 n1303 n785 n210 n815 n829 n845 n859 n875 gng_smul_16_18_sadd_37 
Xu_gng_smul_16_18 SYNOPSYS_UNCONNECTED_4 mul1[32] mul1[31] mul1[30] mul1[29] mul1[28] 
+ mul1[27] mul1[26] mul1[25] mul1[24] mul1[23] mul1[22] mul1[21] mul1[20] mul1[19] 
+ SYNOPSYS_UNCONNECTED_9 SYNOPSYS_UNCONNECTED_8 SYNOPSYS_UNCONNECTED_7 SYNOPSYS_UNCONNECTED_6 
+ SYNOPSYS_UNCONNECTED_5 SYNOPSYS_UNCONNECTED_17 SYNOPSYS_UNCONNECTED_16 SYNOPSYS_UNCONNECTED_15 
+ SYNOPSYS_UNCONNECTED_14 SYNOPSYS_UNCONNECTED_13 SYNOPSYS_UNCONNECTED_12 SYNOPSYS_UNCONNECTED_11 
+ SYNOPSYS_UNCONNECTED_10 SYNOPSYS_UNCONNECTED_23 SYNOPSYS_UNCONNECTED_22 SYNOPSYS_UNCONNECTED_21 
+ SYNOPSYS_UNCONNECTED_20 SYNOPSYS_UNCONNECTED_19 SYNOPSYS_UNCONNECTED_18 n6111 
+ sum1[37] sum1[36] sum1[35] sum1[34] sum1[33] sum1[32] sum1[31] sum1[30] sum1[29] 
+ sum1[28] sum1[27] sum1[26] sum1[25] sum1[24] sum1[23] sum1[22] sum1[21] sum1[20] 
+ VSS n286 n290 n294 n298 n302 n306 n310 n314 n318 n322 n326 n330 n334 n338 n342 gng_smul_16_18 
Xadd_219 N1810 N1800 N1790 N1780 N1770 N1760 N1750 N1740 N1730 N1720 N1710 N1700 
+ N1690 N1680 N1670 SYNOPSYS_UNCONNECTED_3 VDD n29 n30 n31 n32 n33 n34 n35 n36 n37 
+ n38 n39 n40 n41 n42 n43 gng_interp_DW01_inc_0 
Xadd_199 N131 N130 N129 N128 N127 N126 N125 N124 N123 N122 N121 N120 N119 N118 N117 
+ N116 SYNOPSYS_UNCONNECTED_2 SYNOPSYS_UNCONNECTED_1 VSS NETTRAN_DUMMY_16868 mul1[32] 
+ mul1[32] mul1[32] mul1[32] mul1[32] mul1[31] mul1[30] mul1[29] mul1[28] mul1[27] 
+ mul1[26] mul1[25] mul1[24] mul1[23] mul1[22] mul1[21] mul1[20] mul1[19] c0_r5[17] 
+ c0_r5[16] c0_r5[15] c0_r5[14] c0_r5[13] c0_r5[12] c0_r5[11] c0_r5[10] c0_r5[9] 
+ c0_r5[8] c0_r5[7] c0_r5[6] c0_r5[5] c0_r5[4] c0_r5[3] c0_r5[2] c0_r5[1] c0_r5[0] gng_interp_DW01_add_1 
.ENDS

.SUBCKT gng data_out[15] data_out[14] data_out[13] data_out[12] data_out[11] data_out[10] 
+ data_out[9] data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] data_out[3] 
+ data_out[2] data_out[1] data_out[0] valid_out ce rstn clk 
XSPARE_PREFIX_NAME_0_19 VSS VSS NETTRAN_DUMMY_16869 NETTRAN_DUMMY_16870 NETTRAN_DUMMY_16871 NAND2_X4 
XSPARE_PREFIX_NAME_0_18 VSS VSS NETTRAN_DUMMY_16872 NETTRAN_DUMMY_16873 NETTRAN_DUMMY_16874 NAND2_X4 
XSPARE_PREFIX_NAME_0_17 VSS VSS NETTRAN_DUMMY_16875 NETTRAN_DUMMY_16876 NETTRAN_DUMMY_16877 NAND2_X4 
XSPARE_PREFIX_NAME_0_16 VSS VSS NETTRAN_DUMMY_16878 NETTRAN_DUMMY_16879 NETTRAN_DUMMY_16880 NAND2_X4 
XSPARE_PREFIX_NAME_0_15 VSS VSS NETTRAN_DUMMY_16881 NETTRAN_DUMMY_16882 NETTRAN_DUMMY_16883 NAND2_X4 
XSPARE_PREFIX_NAME_0_14 VSS VSS NETTRAN_DUMMY_16884 NETTRAN_DUMMY_16885 NETTRAN_DUMMY_16886 NAND2_X4 
XSPARE_PREFIX_NAME_0_13 VSS VSS NETTRAN_DUMMY_16887 NETTRAN_DUMMY_16888 NETTRAN_DUMMY_16889 NAND2_X4 
XSPARE_PREFIX_NAME_0_12 VSS VSS NETTRAN_DUMMY_16890 NETTRAN_DUMMY_16891 NETTRAN_DUMMY_16892 NAND2_X4 
XSPARE_PREFIX_NAME_0_11 VSS VSS NETTRAN_DUMMY_16893 NETTRAN_DUMMY_16894 NETTRAN_DUMMY_16895 NAND2_X4 
XSPARE_PREFIX_NAME_0_10 VSS VSS NETTRAN_DUMMY_16896 NETTRAN_DUMMY_16897 NETTRAN_DUMMY_16898 NAND2_X4 
XSPARE_PREFIX_NAME_0_9 VSS VSS NETTRAN_DUMMY_16899 NETTRAN_DUMMY_16900 NETTRAN_DUMMY_16901 NAND2_X4 
XSPARE_PREFIX_NAME_0_8 VSS VSS NETTRAN_DUMMY_16902 NETTRAN_DUMMY_16903 NETTRAN_DUMMY_16904 NAND2_X4 
XSPARE_PREFIX_NAME_0_7 VSS VSS NETTRAN_DUMMY_16905 NETTRAN_DUMMY_16906 NETTRAN_DUMMY_16907 NAND2_X4 
XSPARE_PREFIX_NAME_0_6 VSS VSS NETTRAN_DUMMY_16908 NETTRAN_DUMMY_16909 NETTRAN_DUMMY_16910 NAND2_X4 
XSPARE_PREFIX_NAME_0_5 VSS VSS NETTRAN_DUMMY_16911 NETTRAN_DUMMY_16912 NETTRAN_DUMMY_16913 NAND2_X4 
XSPARE_PREFIX_NAME_0_4 VSS VSS NETTRAN_DUMMY_16914 NETTRAN_DUMMY_16915 NETTRAN_DUMMY_16916 NAND2_X4 
XSPARE_PREFIX_NAME_0_3 VSS VSS NETTRAN_DUMMY_16917 NETTRAN_DUMMY_16918 NETTRAN_DUMMY_16919 NAND2_X4 
XSPARE_PREFIX_NAME_0_2 VSS VSS NETTRAN_DUMMY_16920 NETTRAN_DUMMY_16921 NETTRAN_DUMMY_16922 NAND2_X4 
XSPARE_PREFIX_NAME_0_1 VSS VSS NETTRAN_DUMMY_16923 NETTRAN_DUMMY_16924 NETTRAN_DUMMY_16925 NAND2_X4 
XSPARE_PREFIX_NAME_0_0 VSS VSS NETTRAN_DUMMY_16926 NETTRAN_DUMMY_16927 NETTRAN_DUMMY_16928 NAND2_X4 
XSPARE_PREFIX_NAME_19 VSS VSS NETTRAN_DUMMY_16929 NETTRAN_DUMMY_16930 NETTRAN_DUMMY_16931 NOR2_X4 
XSPARE_PREFIX_NAME_18 VSS VSS NETTRAN_DUMMY_16932 NETTRAN_DUMMY_16933 NETTRAN_DUMMY_16934 NOR2_X4 
XSPARE_PREFIX_NAME_17 VSS VSS NETTRAN_DUMMY_16935 NETTRAN_DUMMY_16936 NETTRAN_DUMMY_16937 NOR2_X4 
XSPARE_PREFIX_NAME_16 VSS VSS NETTRAN_DUMMY_16938 NETTRAN_DUMMY_16939 NETTRAN_DUMMY_16940 NOR2_X4 
XSPARE_PREFIX_NAME_15 VSS VSS NETTRAN_DUMMY_16941 NETTRAN_DUMMY_16942 NETTRAN_DUMMY_16943 NOR2_X4 
XSPARE_PREFIX_NAME_14 VSS VSS NETTRAN_DUMMY_16944 NETTRAN_DUMMY_16945 NETTRAN_DUMMY_16946 NOR2_X4 
XSPARE_PREFIX_NAME_13 VSS VSS NETTRAN_DUMMY_16947 NETTRAN_DUMMY_16948 NETTRAN_DUMMY_16949 NOR2_X4 
XSPARE_PREFIX_NAME_12 VSS VSS NETTRAN_DUMMY_16950 NETTRAN_DUMMY_16951 NETTRAN_DUMMY_16952 NOR2_X4 
XSPARE_PREFIX_NAME_11 VSS VSS NETTRAN_DUMMY_16953 NETTRAN_DUMMY_16954 NETTRAN_DUMMY_16955 NOR2_X4 
XSPARE_PREFIX_NAME_10 VSS VSS NETTRAN_DUMMY_16956 NETTRAN_DUMMY_16957 NETTRAN_DUMMY_16958 NOR2_X4 
XSPARE_PREFIX_NAME_9 VSS VSS NETTRAN_DUMMY_16959 NETTRAN_DUMMY_16960 NETTRAN_DUMMY_16961 NOR2_X4 
XSPARE_PREFIX_NAME_8 VSS VSS NETTRAN_DUMMY_16962 NETTRAN_DUMMY_16963 NETTRAN_DUMMY_16964 NOR2_X4 
XSPARE_PREFIX_NAME_7 VSS VSS NETTRAN_DUMMY_16965 NETTRAN_DUMMY_16966 NETTRAN_DUMMY_16967 NOR2_X4 
XSPARE_PREFIX_NAME_6 VSS VSS NETTRAN_DUMMY_16968 NETTRAN_DUMMY_16969 NETTRAN_DUMMY_16970 NOR2_X4 
XSPARE_PREFIX_NAME_5 VSS VSS NETTRAN_DUMMY_16971 NETTRAN_DUMMY_16972 NETTRAN_DUMMY_16973 NOR2_X4 
XSPARE_PREFIX_NAME_4 VSS VSS NETTRAN_DUMMY_16974 NETTRAN_DUMMY_16975 NETTRAN_DUMMY_16976 NOR2_X4 
XSPARE_PREFIX_NAME_3 VSS VSS NETTRAN_DUMMY_16977 NETTRAN_DUMMY_16978 NETTRAN_DUMMY_16979 NOR2_X4 
XSPARE_PREFIX_NAME_2 VSS VSS NETTRAN_DUMMY_16980 NETTRAN_DUMMY_16981 NETTRAN_DUMMY_16982 NOR2_X4 
XSPARE_PREFIX_NAME_1 VSS VSS NETTRAN_DUMMY_16983 NETTRAN_DUMMY_16984 NETTRAN_DUMMY_16985 NOR2_X4 
XSPARE_PREFIX_NAME_0 VSS VSS NETTRAN_DUMMY_16986 NETTRAN_DUMMY_16987 NETTRAN_DUMMY_16988 NOR2_X4 
XU3 rstn n3 NETTRAN_DUMMY_16989 NETTRAN_DUMMY_16990 BUF_X2 
XU2 rstn n2 NETTRAN_DUMMY_16991 NETTRAN_DUMMY_16992 BUF_X1 
XU1 rstn n1 NETTRAN_DUMMY_16993 NETTRAN_DUMMY_16994 BUF_X2 
XCLKBUF_X3_G1B1I9 clk clk_G1B1I9 NETTRAN_DUMMY_16995 NETTRAN_DUMMY_16996 CLKBUF_X1 
Xu_gng_ctg clk n1 ce valid_out_ctg n3 n2 data_out_ctg[63] data_out_ctg[62] data_out_ctg[61] 
+ data_out_ctg[60] data_out_ctg[59] data_out_ctg[58] data_out_ctg[57] data_out_ctg[56] 
+ data_out_ctg[55] data_out_ctg[54] data_out_ctg[53] data_out_ctg[52] data_out_ctg[51] 
+ data_out_ctg[50] data_out_ctg[49] data_out_ctg[48] data_out_ctg[47] data_out_ctg[46] 
+ data_out_ctg[45] data_out_ctg[44] data_out_ctg[43] data_out_ctg[42] data_out_ctg[41] 
+ data_out_ctg[40] data_out_ctg[39] data_out_ctg[38] data_out_ctg[37] data_out_ctg[36] 
+ data_out_ctg[35] data_out_ctg[34] data_out_ctg[33] data_out_ctg[32] data_out_ctg[31] 
+ data_out_ctg[30] data_out_ctg[29] data_out_ctg[28] data_out_ctg[27] data_out_ctg[26] 
+ data_out_ctg[25] data_out_ctg[24] data_out_ctg[23] data_out_ctg[22] data_out_ctg[21] 
+ data_out_ctg[20] data_out_ctg[19] data_out_ctg[18] data_out_ctg[17] data_out_ctg[16] 
+ data_out_ctg[15] data_out_ctg[14] data_out_ctg[13] data_out_ctg[12] data_out_ctg[11] 
+ data_out_ctg[10] data_out_ctg[9] data_out_ctg[8] data_out_ctg[7] data_out_ctg[6] 
+ data_out_ctg[5] data_out_ctg[4] data_out_ctg[3] data_out_ctg[2] data_out_ctg[1] 
+ data_out_ctg[0] n1 rstn clk_G1B1I9 gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff 
Xu_gng_interp clk n2 valid_out_ctg valid_out n3 n2 data_out[15] data_out[14] data_out[13] 
+ data_out[12] data_out[11] data_out[10] data_out[9] data_out[8] data_out[7] data_out[6] 
+ data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] data_out_ctg[63] 
+ data_out_ctg[62] data_out_ctg[61] data_out_ctg[60] data_out_ctg[59] data_out_ctg[58] 
+ data_out_ctg[57] data_out_ctg[56] data_out_ctg[55] data_out_ctg[54] data_out_ctg[53] 
+ data_out_ctg[52] data_out_ctg[51] data_out_ctg[50] data_out_ctg[49] data_out_ctg[48] 
+ data_out_ctg[47] data_out_ctg[46] data_out_ctg[45] data_out_ctg[44] data_out_ctg[43] 
+ data_out_ctg[42] data_out_ctg[41] data_out_ctg[40] data_out_ctg[39] data_out_ctg[38] 
+ data_out_ctg[37] data_out_ctg[36] data_out_ctg[35] data_out_ctg[34] data_out_ctg[33] 
+ data_out_ctg[32] data_out_ctg[31] data_out_ctg[30] data_out_ctg[29] data_out_ctg[28] 
+ data_out_ctg[27] data_out_ctg[26] data_out_ctg[25] data_out_ctg[24] data_out_ctg[23] 
+ data_out_ctg[22] data_out_ctg[21] data_out_ctg[20] data_out_ctg[19] data_out_ctg[18] 
+ data_out_ctg[17] data_out_ctg[16] data_out_ctg[15] data_out_ctg[14] data_out_ctg[13] 
+ data_out_ctg[12] data_out_ctg[11] data_out_ctg[10] data_out_ctg[9] data_out_ctg[8] 
+ data_out_ctg[7] data_out_ctg[6] data_out_ctg[5] data_out_ctg[4] data_out_ctg[3] 
+ data_out_ctg[2] data_out_ctg[1] data_out_ctg[0] n1 clk_G1B1I9 gng_interp 
.ENDS

