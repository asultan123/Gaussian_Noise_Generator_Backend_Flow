
module gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff ( clk, rstn, 
        ce, valid_out, data_out );
  output [63:0] data_out;
  input clk, rstn, ce;
  output valid_out;
  wire   N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n77, n79, n81, n83, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n128, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n2460, n2470, n2480, n2490, n2500, n2510, n2520, n2530,
         n2540, n2550, n2560, n2570, n2580, n2590, n2600, n2610, n2620, n2630,
         n2640, n2650, n2660, n2670, n2680, n2690, n2700, n2710, n2720, n2730,
         n2740, n2750, n2760, n2770, n2780, n2790, n2800, n2810, n2820, n2830,
         n2840, n2850, n2860, n2870, n2880, n2890, n2900, n2910, n2920, n2930,
         n2940, n2950, n2960, n2970, n2980, n2990, n3000, n3010, n3020, n3030,
         n3040, n3050, n3060, n3070, n3080, n3090, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n76, n78, n80, n82, n84,
         n125, n127, n129, n185, n186, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626;
  wire   [54:40] z1;
  wire   [63:25] z1_next;
  wire   [63:61] z2;
  wire   [63:19] z2_next;
  wire   [63:57] z3;
  wire   [63:16] z3_next;

  DFF_X1 z3_reg_9_ ( .D(n551), .CK(clk), .Q(z3_next[16]), .QN(n55) );
  DFF_X1 z3_reg_16_ ( .D(n544), .CK(clk), .Q(z3_next[23]), .QN(n48) );
  DFF_X1 z3_reg_23_ ( .D(n537), .CK(clk), .QN(n41) );
  DFF_X1 z3_reg_30_ ( .D(n530), .CK(clk), .Q(z3_next[37]), .QN(n34) );
  DFF_X1 z3_reg_37_ ( .D(n523), .CK(clk), .Q(z3_next[44]), .QN(n27) );
  DFF_X1 z3_reg_44_ ( .D(n516), .CK(clk), .QN(n20) );
  DFF_X1 z3_reg_51_ ( .D(n509), .CK(clk), .Q(z3_next[58]), .QN(n13) );
  DFF_X1 z3_reg_58_ ( .D(n502), .CK(clk), .Q(z3[58]), .QN(n6) );
  DFF_X1 z3_reg_13_ ( .D(n547), .CK(clk), .Q(z3_next[20]), .QN(n51) );
  DFF_X1 z3_reg_20_ ( .D(n540), .CK(clk), .QN(n44) );
  DFF_X1 z3_reg_27_ ( .D(n533), .CK(clk), .Q(z3_next[34]), .QN(n37) );
  DFF_X1 z3_reg_34_ ( .D(n526), .CK(clk), .Q(z3_next[41]), .QN(n30) );
  DFF_X1 z3_reg_41_ ( .D(n519), .CK(clk), .QN(n23) );
  DFF_X1 z3_reg_48_ ( .D(n512), .CK(clk), .QN(n16) );
  DFF_X1 z3_reg_55_ ( .D(n505), .CK(clk), .Q(z3_next[62]), .QN(n9) );
  DFF_X1 z3_reg_62_ ( .D(n498), .CK(clk), .Q(z3[62]), .QN(n2) );
  DFF_X1 z3_reg_10_ ( .D(n550), .CK(clk), .Q(z3_next[17]), .QN(n54) );
  DFF_X1 z3_reg_17_ ( .D(n543), .CK(clk), .Q(z3_next[24]), .QN(n47) );
  DFF_X1 z3_reg_24_ ( .D(n536), .CK(clk), .Q(z3_next[31]), .QN(n40) );
  DFF_X1 z3_reg_31_ ( .D(n529), .CK(clk), .Q(z3_next[38]), .QN(n33) );
  DFF_X1 z3_reg_38_ ( .D(n522), .CK(clk), .Q(z3_next[45]), .QN(n26) );
  DFF_X1 z3_reg_45_ ( .D(n515), .CK(clk), .QN(n19) );
  DFF_X1 z3_reg_52_ ( .D(n508), .CK(clk), .QN(n12) );
  DFF_X1 z3_reg_59_ ( .D(n501), .CK(clk), .Q(z3[59]), .QN(n5) );
  DFF_X1 z3_reg_14_ ( .D(n546), .CK(clk), .Q(z3_next[21]), .QN(n50) );
  DFF_X1 z3_reg_21_ ( .D(n539), .CK(clk), .QN(n43) );
  DFF_X1 z3_reg_28_ ( .D(n532), .CK(clk), .Q(z3_next[35]), .QN(n36) );
  DFF_X1 z3_reg_35_ ( .D(n525), .CK(clk), .Q(z3_next[42]), .QN(n29) );
  DFF_X1 z3_reg_42_ ( .D(n518), .CK(clk), .QN(n22) );
  DFF_X1 z3_reg_49_ ( .D(n511), .CK(clk), .QN(n15) );
  DFF_X1 z3_reg_56_ ( .D(n504), .CK(clk), .Q(z3_next[63]), .QN(n8) );
  DFF_X1 z3_reg_63_ ( .D(n497), .CK(clk), .Q(z3[63]), .QN(n1) );
  DFF_X1 z3_reg_11_ ( .D(n549), .CK(clk), .Q(z3_next[18]), .QN(n53) );
  DFF_X1 z3_reg_18_ ( .D(n542), .CK(clk), .QN(n46) );
  DFF_X1 z3_reg_25_ ( .D(n535), .CK(clk), .Q(z3_next[32]), .QN(n39) );
  DFF_X1 z3_reg_32_ ( .D(n528), .CK(clk), .Q(z3_next[39]), .QN(n32) );
  DFF_X1 z3_reg_39_ ( .D(n521), .CK(clk), .Q(z3_next[46]), .QN(n25) );
  DFF_X1 z3_reg_46_ ( .D(n514), .CK(clk), .QN(n18) );
  DFF_X1 z3_reg_53_ ( .D(n507), .CK(clk), .QN(n11) );
  DFF_X1 z3_reg_60_ ( .D(n500), .CK(clk), .Q(z3[60]), .QN(n4) );
  DFF_X1 z3_reg_15_ ( .D(n545), .CK(clk), .Q(z3_next[22]), .QN(n49) );
  DFF_X1 z3_reg_22_ ( .D(n538), .CK(clk), .QN(n42) );
  DFF_X1 z3_reg_29_ ( .D(n531), .CK(clk), .Q(z3_next[36]), .QN(n35) );
  DFF_X1 z3_reg_36_ ( .D(n524), .CK(clk), .Q(z3_next[43]), .QN(n28) );
  DFF_X1 z3_reg_43_ ( .D(n517), .CK(clk), .QN(n21) );
  DFF_X1 z3_reg_50_ ( .D(n510), .CK(clk), .QN(n14) );
  DFF_X1 z3_reg_57_ ( .D(n503), .CK(clk), .Q(z3[57]), .QN(n7) );
  DFF_X1 z3_reg_12_ ( .D(n548), .CK(clk), .Q(z3_next[19]), .QN(n52) );
  DFF_X1 z3_reg_19_ ( .D(n541), .CK(clk), .QN(n45) );
  DFF_X1 z3_reg_26_ ( .D(n534), .CK(clk), .Q(z3_next[33]), .QN(n38) );
  DFF_X1 z3_reg_33_ ( .D(n527), .CK(clk), .Q(z3_next[40]), .QN(n31) );
  DFF_X1 z3_reg_40_ ( .D(n520), .CK(clk), .QN(n24) );
  DFF_X1 z3_reg_47_ ( .D(n513), .CK(clk), .QN(n17) );
  DFF_X1 z3_reg_54_ ( .D(n506), .CK(clk), .Q(z3_next[61]), .QN(n10) );
  DFF_X1 z3_reg_61_ ( .D(n499), .CK(clk), .Q(z3[61]), .QN(n3) );
  DFF_X1 z1_reg_1_ ( .D(n496), .CK(clk), .Q(z1_next[25]), .QN(n123) );
  DFF_X1 z1_reg_25_ ( .D(n472), .CK(clk), .Q(z1_next[49]), .QN(n99) );
  DFF_X1 z1_reg_49_ ( .D(n448), .CK(clk), .Q(z1[49]), .QN(n70) );
  DFF_X1 z1_reg_15_ ( .D(n482), .CK(clk), .Q(z1_next[39]), .QN(n109) );
  DFF_X1 z1_reg_39_ ( .D(n458), .CK(clk), .Q(z1_next[63]), .QN(n85) );
  DFF_X1 z1_reg_63_ ( .D(n434), .CK(clk), .QN(n56) );
  DFF_X1 z1_reg_5_ ( .D(n492), .CK(clk), .Q(z1_next[29]), .QN(n119) );
  DFF_X1 z1_reg_29_ ( .D(n468), .CK(clk), .Q(z1_next[53]), .QN(n95) );
  DFF_X1 z1_reg_53_ ( .D(n444), .CK(clk), .Q(z1[53]), .QN(n66) );
  DFF_X1 z1_reg_19_ ( .D(n478), .CK(clk), .Q(z1_next[43]), .QN(n105) );
  DFF_X1 z1_reg_43_ ( .D(n454), .CK(clk), .Q(z1[43]), .QN(n77) );
  DFF_X1 z1_reg_4_ ( .D(n493), .CK(clk), .Q(z1_next[28]), .QN(n120) );
  DFF_X1 z1_reg_28_ ( .D(n469), .CK(clk), .Q(z1_next[52]), .QN(n96) );
  DFF_X1 z1_reg_52_ ( .D(n445), .CK(clk), .Q(z1[52]), .QN(n67) );
  DFF_X1 z1_reg_18_ ( .D(n479), .CK(clk), .Q(z1_next[42]), .QN(n106) );
  DFF_X1 z1_reg_42_ ( .D(n455), .CK(clk), .Q(z1[42]), .QN(n79) );
  DFF_X1 z1_reg_3_ ( .D(n494), .CK(clk), .Q(z1_next[27]), .QN(n121) );
  DFF_X1 z1_reg_27_ ( .D(n470), .CK(clk), .Q(z1_next[51]), .QN(n97) );
  DFF_X1 z1_reg_51_ ( .D(n446), .CK(clk), .Q(z1[51]), .QN(n68) );
  DFF_X1 z1_reg_17_ ( .D(n480), .CK(clk), .Q(z1_next[41]), .QN(n107) );
  DFF_X1 z1_reg_41_ ( .D(n456), .CK(clk), .Q(z1[41]), .QN(n81) );
  DFF_X1 z1_reg_2_ ( .D(n495), .CK(clk), .Q(z1_next[26]), .QN(n122) );
  DFF_X1 z1_reg_26_ ( .D(n471), .CK(clk), .Q(z1_next[50]), .QN(n98) );
  DFF_X1 z1_reg_50_ ( .D(n447), .CK(clk), .Q(z1[50]), .QN(n69) );
  DFF_X1 z1_reg_16_ ( .D(n481), .CK(clk), .Q(z1_next[40]), .QN(n108) );
  DFF_X1 z1_reg_40_ ( .D(n457), .CK(clk), .Q(z1[40]), .QN(n83) );
  DFF_X1 z1_reg_6_ ( .D(n491), .CK(clk), .Q(z1_next[30]), .QN(n118) );
  DFF_X1 z1_reg_30_ ( .D(n467), .CK(clk), .Q(z1_next[54]), .QN(n94) );
  DFF_X1 z1_reg_54_ ( .D(n443), .CK(clk), .Q(z1[54]), .QN(n65) );
  DFF_X1 z1_reg_20_ ( .D(n477), .CK(clk), .Q(z1_next[44]), .QN(n104) );
  DFF_X1 z1_reg_44_ ( .D(n453), .CK(clk), .Q(z1[44]), .QN(n75) );
  DFF_X1 z1_reg_10_ ( .D(n487), .CK(clk), .Q(z1_next[34]), .QN(n114) );
  DFF_X1 z1_reg_34_ ( .D(n463), .CK(clk), .QN(n90) );
  DFF_X1 z1_reg_58_ ( .D(n439), .CK(clk), .QN(n61) );
  DFF_X1 z1_reg_24_ ( .D(n473), .CK(clk), .Q(z1_next[48]), .QN(n100) );
  DFF_X1 z1_reg_48_ ( .D(n449), .CK(clk), .Q(z1[48]), .QN(n71) );
  DFF_X1 z1_reg_9_ ( .D(n488), .CK(clk), .Q(z1_next[33]), .QN(n115) );
  DFF_X1 z1_reg_33_ ( .D(n464), .CK(clk), .Q(z1_next[57]), .QN(n91) );
  DFF_X1 z1_reg_57_ ( .D(n440), .CK(clk), .QN(n62) );
  DFF_X1 z1_reg_14_ ( .D(n483), .CK(clk), .Q(z1_next[38]), .QN(n110) );
  DFF_X1 z1_reg_38_ ( .D(n459), .CK(clk), .Q(z1_next[62]), .QN(n86) );
  DFF_X1 z1_reg_62_ ( .D(n435), .CK(clk), .QN(n57) );
  DFF_X1 z1_reg_23_ ( .D(n474), .CK(clk), .Q(z1_next[47]), .QN(n101) );
  DFF_X1 z1_reg_47_ ( .D(n450), .CK(clk), .Q(z1[47]), .QN(n72) );
  DFF_X1 z1_reg_8_ ( .D(n489), .CK(clk), .Q(z1_next[32]), .QN(n116) );
  DFF_X1 z1_reg_32_ ( .D(n465), .CK(clk), .Q(z1_next[56]), .QN(n92) );
  DFF_X1 z1_reg_56_ ( .D(n441), .CK(clk), .QN(n63) );
  DFF_X1 z1_reg_13_ ( .D(n484), .CK(clk), .Q(z1_next[37]), .QN(n111) );
  DFF_X1 z1_reg_37_ ( .D(n460), .CK(clk), .Q(z1_next[61]), .QN(n87) );
  DFF_X1 z1_reg_61_ ( .D(n436), .CK(clk), .QN(n58) );
  DFF_X1 z1_reg_22_ ( .D(n475), .CK(clk), .Q(z1_next[46]), .QN(n102) );
  DFF_X1 z1_reg_46_ ( .D(n451), .CK(clk), .Q(z1[46]), .QN(n73) );
  DFF_X1 z1_reg_7_ ( .D(n490), .CK(clk), .Q(z1_next[31]), .QN(n117) );
  DFF_X1 z1_reg_31_ ( .D(n466), .CK(clk), .Q(z1_next[55]), .QN(n93) );
  DFF_X1 z1_reg_55_ ( .D(n442), .CK(clk), .QN(n64) );
  DFF_X1 z1_reg_12_ ( .D(n485), .CK(clk), .Q(z1_next[36]), .QN(n112) );
  DFF_X1 z1_reg_36_ ( .D(n461), .CK(clk), .Q(z1_next[60]), .QN(n88) );
  DFF_X1 z1_reg_60_ ( .D(n437), .CK(clk), .QN(n59) );
  DFF_X1 z1_reg_21_ ( .D(n476), .CK(clk), .Q(z1_next[45]), .QN(n103) );
  DFF_X1 z1_reg_45_ ( .D(n452), .CK(clk), .Q(z1[45]), .QN(n74) );
  DFF_X1 z1_reg_11_ ( .D(n486), .CK(clk), .Q(z1_next[35]), .QN(n113) );
  DFF_X1 z1_reg_35_ ( .D(n462), .CK(clk), .Q(z1_next[59]), .QN(n89) );
  DFF_X1 z1_reg_59_ ( .D(n438), .CK(clk), .QN(n60) );
  DFF_X1 z2_reg_6_ ( .D(n433), .CK(clk), .Q(z2_next[19]), .QN(n184) );
  DFF_X1 z2_reg_19_ ( .D(n420), .CK(clk), .Q(z2_next[32]), .QN(n171) );
  DFF_X1 z2_reg_32_ ( .D(n407), .CK(clk), .Q(z2_next[45]), .QN(n158) );
  DFF_X1 z2_reg_45_ ( .D(n394), .CK(clk), .Q(z2_next[58]), .QN(n145) );
  DFF_X1 z2_reg_58_ ( .D(n381), .CK(clk), .QN(n132) );
  DFF_X1 z2_reg_13_ ( .D(n426), .CK(clk), .Q(z2_next[26]), .QN(n177) );
  DFF_X1 z2_reg_26_ ( .D(n413), .CK(clk), .Q(z2_next[39]), .QN(n164) );
  DFF_X1 z2_reg_39_ ( .D(n400), .CK(clk), .Q(z2_next[52]), .QN(n151) );
  DFF_X1 z2_reg_52_ ( .D(n387), .CK(clk), .QN(n138) );
  DFF_X1 z2_reg_7_ ( .D(n432), .CK(clk), .Q(z2_next[20]), .QN(n183) );
  DFF_X1 z2_reg_20_ ( .D(n419), .CK(clk), .Q(z2_next[33]), .QN(n170) );
  DFF_X1 z2_reg_33_ ( .D(n406), .CK(clk), .Q(z2_next[46]), .QN(n157) );
  DFF_X1 z2_reg_46_ ( .D(n393), .CK(clk), .Q(z2_next[59]), .QN(n144) );
  DFF_X1 z2_reg_59_ ( .D(n380), .CK(clk), .QN(n131) );
  DFF_X1 z2_reg_14_ ( .D(n425), .CK(clk), .Q(z2_next[27]), .QN(n176) );
  DFF_X1 z2_reg_27_ ( .D(n412), .CK(clk), .Q(z2_next[40]), .QN(n163) );
  DFF_X1 z2_reg_40_ ( .D(n399), .CK(clk), .Q(z2_next[53]), .QN(n150) );
  DFF_X1 z2_reg_53_ ( .D(n386), .CK(clk), .QN(n137) );
  DFF_X1 z2_reg_8_ ( .D(n431), .CK(clk), .Q(z2_next[21]), .QN(n182) );
  DFF_X1 z2_reg_21_ ( .D(n418), .CK(clk), .Q(z2_next[34]), .QN(n169) );
  DFF_X1 z2_reg_34_ ( .D(n405), .CK(clk), .Q(z2_next[47]), .QN(n156) );
  DFF_X1 z2_reg_47_ ( .D(n392), .CK(clk), .Q(z2_next[60]), .QN(n143) );
  DFF_X1 z2_reg_60_ ( .D(n379), .CK(clk), .QN(n130) );
  DFF_X1 z2_reg_15_ ( .D(n424), .CK(clk), .Q(z2_next[28]), .QN(n175) );
  DFF_X1 z2_reg_28_ ( .D(n411), .CK(clk), .Q(z2_next[41]), .QN(n162) );
  DFF_X1 z2_reg_41_ ( .D(n398), .CK(clk), .Q(z2_next[54]), .QN(n149) );
  DFF_X1 z2_reg_54_ ( .D(n385), .CK(clk), .QN(n136) );
  DFF_X1 z2_reg_9_ ( .D(n430), .CK(clk), .Q(z2_next[22]), .QN(n181) );
  DFF_X1 z2_reg_22_ ( .D(n417), .CK(clk), .Q(z2_next[35]), .QN(n168) );
  DFF_X1 z2_reg_35_ ( .D(n404), .CK(clk), .Q(z2_next[48]), .QN(n155) );
  DFF_X1 z2_reg_48_ ( .D(n391), .CK(clk), .Q(z2_next[61]), .QN(n142) );
  DFF_X1 z2_reg_61_ ( .D(n378), .CK(clk), .Q(z2[61]), .QN(n128) );
  DFF_X1 z2_reg_16_ ( .D(n423), .CK(clk), .Q(z2_next[29]), .QN(n174) );
  DFF_X1 z2_reg_29_ ( .D(n410), .CK(clk), .Q(z2_next[42]), .QN(n161) );
  DFF_X1 z2_reg_42_ ( .D(n397), .CK(clk), .Q(z2_next[55]), .QN(n148) );
  DFF_X1 z2_reg_55_ ( .D(n384), .CK(clk), .QN(n135) );
  DFF_X1 z2_reg_10_ ( .D(n429), .CK(clk), .Q(z2_next[23]), .QN(n180) );
  DFF_X1 z2_reg_23_ ( .D(n416), .CK(clk), .Q(z2_next[36]), .QN(n167) );
  DFF_X1 z2_reg_36_ ( .D(n403), .CK(clk), .Q(z2_next[49]), .QN(n154) );
  DFF_X1 z2_reg_49_ ( .D(n390), .CK(clk), .Q(z2_next[62]), .QN(n141) );
  DFF_X1 z2_reg_62_ ( .D(n377), .CK(clk), .Q(z2[62]), .QN(n126) );
  DFF_X1 z2_reg_17_ ( .D(n422), .CK(clk), .Q(z2_next[30]), .QN(n173) );
  DFF_X1 z2_reg_30_ ( .D(n409), .CK(clk), .Q(z2_next[43]), .QN(n160) );
  DFF_X1 z2_reg_43_ ( .D(n396), .CK(clk), .Q(z2_next[56]), .QN(n147) );
  DFF_X1 z2_reg_56_ ( .D(n383), .CK(clk), .QN(n134) );
  DFF_X1 z2_reg_11_ ( .D(n428), .CK(clk), .Q(z2_next[24]), .QN(n179) );
  DFF_X1 z2_reg_24_ ( .D(n415), .CK(clk), .Q(z2_next[37]), .QN(n166) );
  DFF_X1 z2_reg_37_ ( .D(n402), .CK(clk), .Q(z2_next[50]), .QN(n153) );
  DFF_X1 z2_reg_50_ ( .D(n389), .CK(clk), .Q(z2_next[63]), .QN(n140) );
  DFF_X1 z2_reg_63_ ( .D(n376), .CK(clk), .Q(z2[63]), .QN(n124) );
  DFF_X1 z2_reg_18_ ( .D(n421), .CK(clk), .Q(z2_next[31]), .QN(n172) );
  DFF_X1 z2_reg_31_ ( .D(n408), .CK(clk), .Q(z2_next[44]), .QN(n159) );
  DFF_X1 z2_reg_44_ ( .D(n395), .CK(clk), .Q(z2_next[57]), .QN(n146) );
  DFF_X1 z2_reg_57_ ( .D(n382), .CK(clk), .QN(n133) );
  DFF_X1 z2_reg_12_ ( .D(n427), .CK(clk), .Q(z2_next[25]), .QN(n178) );
  DFF_X1 z2_reg_25_ ( .D(n414), .CK(clk), .Q(z2_next[38]), .QN(n165) );
  DFF_X1 z2_reg_38_ ( .D(n401), .CK(clk), .Q(z2_next[51]), .QN(n152) );
  DFF_X1 z2_reg_51_ ( .D(n388), .CK(clk), .QN(n139) );
  DFF_X1 valid_out_reg ( .D(n568), .CK(clk), .Q(valid_out) );
  DFF_X1 data_out_reg_63_ ( .D(N309), .CK(clk), .Q(data_out[63]) );
  DFF_X1 data_out_reg_62_ ( .D(N308), .CK(clk), .Q(data_out[62]) );
  DFF_X1 data_out_reg_61_ ( .D(N307), .CK(clk), .Q(data_out[61]) );
  DFF_X1 data_out_reg_60_ ( .D(N306), .CK(clk), .Q(data_out[60]) );
  DFF_X1 data_out_reg_59_ ( .D(N305), .CK(clk), .Q(data_out[59]) );
  DFF_X1 data_out_reg_58_ ( .D(N304), .CK(clk), .Q(data_out[58]) );
  DFF_X1 data_out_reg_57_ ( .D(N303), .CK(clk), .Q(data_out[57]) );
  DFF_X1 data_out_reg_56_ ( .D(N302), .CK(clk), .Q(data_out[56]) );
  DFF_X1 data_out_reg_55_ ( .D(N301), .CK(clk), .Q(data_out[55]) );
  DFF_X1 data_out_reg_54_ ( .D(N300), .CK(clk), .Q(data_out[54]) );
  DFF_X1 data_out_reg_53_ ( .D(N299), .CK(clk), .Q(data_out[53]) );
  DFF_X1 data_out_reg_52_ ( .D(N298), .CK(clk), .Q(data_out[52]) );
  DFF_X1 data_out_reg_51_ ( .D(N297), .CK(clk), .Q(data_out[51]) );
  DFF_X1 data_out_reg_50_ ( .D(N296), .CK(clk), .Q(data_out[50]) );
  DFF_X1 data_out_reg_49_ ( .D(N295), .CK(clk), .Q(data_out[49]) );
  DFF_X1 data_out_reg_48_ ( .D(N294), .CK(clk), .Q(data_out[48]) );
  DFF_X1 data_out_reg_47_ ( .D(N293), .CK(clk), .Q(data_out[47]) );
  DFF_X1 data_out_reg_46_ ( .D(N292), .CK(clk), .Q(data_out[46]) );
  DFF_X1 data_out_reg_45_ ( .D(N291), .CK(clk), .Q(data_out[45]) );
  DFF_X1 data_out_reg_44_ ( .D(N290), .CK(clk), .Q(data_out[44]) );
  DFF_X1 data_out_reg_43_ ( .D(N289), .CK(clk), .Q(data_out[43]) );
  DFF_X1 data_out_reg_42_ ( .D(N288), .CK(clk), .Q(data_out[42]) );
  DFF_X1 data_out_reg_41_ ( .D(N287), .CK(clk), .Q(data_out[41]) );
  DFF_X1 data_out_reg_40_ ( .D(N286), .CK(clk), .Q(data_out[40]) );
  DFF_X1 data_out_reg_39_ ( .D(N285), .CK(clk), .Q(data_out[39]) );
  DFF_X1 data_out_reg_38_ ( .D(N284), .CK(clk), .Q(data_out[38]) );
  DFF_X1 data_out_reg_37_ ( .D(N283), .CK(clk), .Q(data_out[37]) );
  DFF_X1 data_out_reg_36_ ( .D(N282), .CK(clk), .Q(data_out[36]) );
  DFF_X1 data_out_reg_35_ ( .D(N281), .CK(clk), .Q(data_out[35]) );
  DFF_X1 data_out_reg_34_ ( .D(N280), .CK(clk), .Q(data_out[34]) );
  DFF_X1 data_out_reg_33_ ( .D(N279), .CK(clk), .Q(data_out[33]) );
  DFF_X1 data_out_reg_32_ ( .D(N278), .CK(clk), .Q(data_out[32]) );
  DFF_X1 data_out_reg_31_ ( .D(N277), .CK(clk), .Q(data_out[31]) );
  DFF_X1 data_out_reg_30_ ( .D(N276), .CK(clk), .Q(data_out[30]) );
  DFF_X1 data_out_reg_29_ ( .D(N275), .CK(clk), .Q(data_out[29]) );
  DFF_X1 data_out_reg_28_ ( .D(N274), .CK(clk), .Q(data_out[28]) );
  DFF_X1 data_out_reg_27_ ( .D(N273), .CK(clk), .Q(data_out[27]) );
  DFF_X1 data_out_reg_26_ ( .D(N272), .CK(clk), .Q(data_out[26]) );
  DFF_X1 data_out_reg_25_ ( .D(N271), .CK(clk), .Q(data_out[25]) );
  DFF_X1 data_out_reg_24_ ( .D(N270), .CK(clk), .Q(data_out[24]) );
  DFF_X1 data_out_reg_23_ ( .D(N269), .CK(clk), .Q(data_out[23]) );
  DFF_X1 data_out_reg_22_ ( .D(N268), .CK(clk), .Q(data_out[22]) );
  DFF_X1 data_out_reg_21_ ( .D(N267), .CK(clk), .Q(data_out[21]) );
  DFF_X1 data_out_reg_20_ ( .D(N266), .CK(clk), .Q(data_out[20]) );
  DFF_X1 data_out_reg_19_ ( .D(N265), .CK(clk), .Q(data_out[19]) );
  DFF_X1 data_out_reg_18_ ( .D(N264), .CK(clk), .Q(data_out[18]) );
  DFF_X1 data_out_reg_17_ ( .D(N263), .CK(clk), .Q(data_out[17]) );
  DFF_X1 data_out_reg_16_ ( .D(N262), .CK(clk), .Q(data_out[16]) );
  DFF_X1 data_out_reg_15_ ( .D(N261), .CK(clk), .Q(data_out[15]) );
  DFF_X1 data_out_reg_14_ ( .D(N260), .CK(clk), .Q(data_out[14]) );
  DFF_X1 data_out_reg_13_ ( .D(N259), .CK(clk), .Q(data_out[13]) );
  DFF_X1 data_out_reg_12_ ( .D(N258), .CK(clk), .Q(data_out[12]) );
  DFF_X1 data_out_reg_11_ ( .D(N257), .CK(clk), .Q(data_out[11]) );
  DFF_X1 data_out_reg_10_ ( .D(N256), .CK(clk), .Q(data_out[10]) );
  DFF_X1 data_out_reg_9_ ( .D(N255), .CK(clk), .Q(data_out[9]) );
  DFF_X1 data_out_reg_8_ ( .D(N254), .CK(clk), .Q(data_out[8]) );
  DFF_X1 data_out_reg_7_ ( .D(N253), .CK(clk), .Q(data_out[7]) );
  DFF_X1 data_out_reg_6_ ( .D(N252), .CK(clk), .Q(data_out[6]) );
  DFF_X1 data_out_reg_5_ ( .D(N251), .CK(clk), .Q(data_out[5]) );
  DFF_X1 data_out_reg_4_ ( .D(N250), .CK(clk), .Q(data_out[4]) );
  DFF_X1 data_out_reg_3_ ( .D(N249), .CK(clk), .Q(data_out[3]) );
  DFF_X1 data_out_reg_2_ ( .D(N248), .CK(clk), .Q(data_out[2]) );
  DFF_X1 data_out_reg_1_ ( .D(N247), .CK(clk), .Q(data_out[1]) );
  DFF_X1 data_out_reg_0_ ( .D(N246), .CK(clk), .Q(data_out[0]) );
  XOR2_X1 U406 ( .A(n226), .B(n330), .Z(n329) );
  XOR2_X1 U407 ( .A(n192), .B(n211), .Z(n330) );
  XOR2_X1 U408 ( .A(n70), .B(z1[54]), .Z(n211) );
  XOR2_X1 U409 ( .A(n227), .B(n332), .Z(n331) );
  XOR2_X1 U410 ( .A(n193), .B(n212), .Z(n332) );
  XOR2_X1 U411 ( .A(n71), .B(z1[53]), .Z(n212) );
  XOR2_X1 U412 ( .A(n228), .B(n334), .Z(n333) );
  XOR2_X1 U413 ( .A(n194), .B(n213), .Z(n334) );
  XOR2_X1 U414 ( .A(n72), .B(z1[52]), .Z(n213) );
  XOR2_X1 U415 ( .A(n229), .B(n336), .Z(n335) );
  XOR2_X1 U416 ( .A(n195), .B(n214), .Z(n336) );
  XOR2_X1 U417 ( .A(n73), .B(z1[51]), .Z(n214) );
  XOR2_X1 U418 ( .A(n230), .B(n338), .Z(n337) );
  XOR2_X1 U419 ( .A(n196), .B(n215), .Z(n338) );
  XOR2_X1 U420 ( .A(n74), .B(z1[50]), .Z(n215) );
  XOR2_X1 U421 ( .A(n231), .B(n340), .Z(n339) );
  XOR2_X1 U422 ( .A(n197), .B(n216), .Z(n340) );
  XOR2_X1 U423 ( .A(n75), .B(z1[49]), .Z(n216) );
  XOR2_X1 U424 ( .A(n232), .B(n342), .Z(n341) );
  XOR2_X1 U425 ( .A(n198), .B(n217), .Z(n342) );
  XOR2_X1 U426 ( .A(n77), .B(z1[48]), .Z(n217) );
  XOR2_X1 U427 ( .A(n344), .B(n345), .Z(n343) );
  XOR2_X1 U428 ( .A(n199), .B(n218), .Z(n345) );
  XOR2_X1 U429 ( .A(n79), .B(z1[47]), .Z(n218) );
  XOR2_X1 U430 ( .A(n347), .B(n348), .Z(n346) );
  XOR2_X1 U431 ( .A(n200), .B(n219), .Z(n348) );
  XOR2_X1 U432 ( .A(n81), .B(z1[46]), .Z(n219) );
  XOR2_X1 U433 ( .A(n350), .B(n351), .Z(n349) );
  XOR2_X1 U434 ( .A(n201), .B(n220), .Z(n351) );
  XOR2_X1 U435 ( .A(n83), .B(z1[45]), .Z(n220) );
  XOR2_X1 U436 ( .A(n353), .B(n354), .Z(n352) );
  XOR2_X1 U437 ( .A(n357), .B(n358), .Z(n356) );
  XOR2_X1 U438 ( .A(n361), .B(n362), .Z(n360) );
  XOR2_X1 U439 ( .A(n365), .B(n366), .Z(n364) );
  XOR2_X1 U440 ( .A(n369), .B(n370), .Z(n368) );
  XOR2_X1 U441 ( .A(n373), .B(n374), .Z(n372) );
  BUF_X1 U3 ( .A(n76), .Z(n84) );
  BUF_X1 U4 ( .A(n76), .Z(n125) );
  BUF_X1 U5 ( .A(n76), .Z(n127) );
  BUF_X1 U6 ( .A(n76), .Z(n129) );
  BUF_X1 U7 ( .A(n78), .Z(n185) );
  BUF_X1 U8 ( .A(n78), .Z(n186) );
  BUF_X1 U9 ( .A(n78), .Z(n552) );
  BUF_X1 U10 ( .A(n78), .Z(n554) );
  BUF_X1 U11 ( .A(n80), .Z(n555) );
  BUF_X1 U12 ( .A(n78), .Z(n553) );
  BUF_X1 U13 ( .A(n80), .Z(n556) );
  BUF_X1 U14 ( .A(n80), .Z(n557) );
  BUF_X1 U15 ( .A(n76), .Z(n82) );
  BUF_X1 U16 ( .A(n188), .Z(n78) );
  BUF_X1 U17 ( .A(n188), .Z(n76) );
  BUF_X1 U18 ( .A(n188), .Z(n80) );
  NAND2_X1 U19 ( .A1(n578), .A2(n187), .ZN(n188) );
  INV_X1 U20 ( .A(n611), .ZN(n570) );
  INV_X1 U21 ( .A(n611), .ZN(n571) );
  INV_X1 U22 ( .A(n611), .ZN(n572) );
  INV_X1 U23 ( .A(n612), .ZN(n573) );
  INV_X1 U24 ( .A(n612), .ZN(n574) );
  INV_X1 U25 ( .A(n612), .ZN(n575) );
  INV_X1 U26 ( .A(n613), .ZN(n576) );
  INV_X1 U27 ( .A(n613), .ZN(n577) );
  INV_X1 U28 ( .A(n568), .ZN(n559) );
  INV_X1 U29 ( .A(n568), .ZN(n560) );
  INV_X1 U30 ( .A(n187), .ZN(n568) );
  NOR2_X1 U31 ( .A1(n606), .A2(n341), .ZN(N255) );
  NOR2_X1 U32 ( .A1(n605), .A2(n339), .ZN(N256) );
  NOR2_X1 U33 ( .A1(n605), .A2(n337), .ZN(N257) );
  NOR2_X1 U34 ( .A1(n604), .A2(n335), .ZN(N258) );
  NOR2_X1 U35 ( .A1(n604), .A2(n333), .ZN(N259) );
  NOR2_X1 U36 ( .A1(n603), .A2(n331), .ZN(N260) );
  NOR2_X1 U37 ( .A1(n603), .A2(n329), .ZN(N261) );
  OAI221_X1 U38 ( .B1(n561), .B2(n140), .C1(n553), .C2(n124), .A(n574), .ZN(
        n376) );
  OAI221_X1 U39 ( .B1(n561), .B2(n113), .C1(n554), .C2(n89), .A(n573), .ZN(
        n462) );
  OAI221_X1 U40 ( .B1(n561), .B2(n112), .C1(n554), .C2(n88), .A(n573), .ZN(
        n461) );
  OAI221_X1 U41 ( .B1(n561), .B2(n117), .C1(n555), .C2(n93), .A(n574), .ZN(
        n466) );
  OAI221_X1 U42 ( .B1(n561), .B2(n111), .C1(n554), .C2(n87), .A(n573), .ZN(
        n460) );
  OAI221_X1 U43 ( .B1(n561), .B2(n116), .C1(n554), .C2(n92), .A(n574), .ZN(
        n465) );
  OAI221_X1 U44 ( .B1(n561), .B2(n110), .C1(n554), .C2(n86), .A(n573), .ZN(
        n459) );
  OAI221_X1 U45 ( .B1(n562), .B2(n115), .C1(n554), .C2(n91), .A(n573), .ZN(
        n464) );
  OAI221_X1 U46 ( .B1(n561), .B2(n114), .C1(n554), .C2(n90), .A(n573), .ZN(
        n463) );
  OAI221_X1 U47 ( .B1(n561), .B2(n94), .C1(n554), .C2(n65), .A(n573), .ZN(n443) );
  OAI221_X1 U48 ( .B1(n561), .B2(n118), .C1(n555), .C2(n94), .A(n574), .ZN(
        n467) );
  OAI221_X1 U49 ( .B1(n562), .B2(n122), .C1(n555), .C2(n98), .A(n574), .ZN(
        n471) );
  OAI221_X1 U50 ( .B1(n562), .B2(n121), .C1(n555), .C2(n97), .A(n574), .ZN(
        n470) );
  OAI221_X1 U51 ( .B1(n561), .B2(n96), .C1(n554), .C2(n67), .A(n573), .ZN(n445) );
  OAI221_X1 U52 ( .B1(n562), .B2(n120), .C1(n555), .C2(n96), .A(n574), .ZN(
        n469) );
  OAI221_X1 U53 ( .B1(n562), .B2(n119), .C1(n555), .C2(n95), .A(n574), .ZN(
        n468) );
  OAI221_X1 U54 ( .B1(n561), .B2(n109), .C1(n554), .C2(n85), .A(n573), .ZN(
        n458) );
  OAI221_X1 U55 ( .B1(n562), .B2(n123), .C1(n555), .C2(n99), .A(n574), .ZN(
        n472) );
  OAI221_X1 U56 ( .B1(n563), .B2(n10), .C1(n556), .C2(n3), .A(n576), .ZN(n499)
         );
  OAI221_X1 U57 ( .B1(n563), .B2(n17), .C1(n557), .C2(n10), .A(n576), .ZN(n506) );
  OAI221_X1 U58 ( .B1(n562), .B2(n52), .C1(n558), .C2(n45), .A(n577), .ZN(n541) );
  OAI221_X1 U59 ( .B1(n563), .B2(n14), .C1(n557), .C2(n7), .A(n576), .ZN(n503)
         );
  OAI221_X1 U60 ( .B1(n563), .B2(n49), .C1(n558), .C2(n42), .A(n577), .ZN(n538) );
  OAI221_X1 U61 ( .B1(n562), .B2(n11), .C1(n556), .C2(n4), .A(n576), .ZN(n500)
         );
  OAI221_X1 U62 ( .B1(n562), .B2(n8), .C1(n556), .C2(n1), .A(n575), .ZN(n497)
         );
  OAI221_X1 U63 ( .B1(n562), .B2(n15), .C1(n557), .C2(n8), .A(n576), .ZN(n504)
         );
  OAI221_X1 U64 ( .B1(n563), .B2(n22), .C1(n557), .C2(n15), .A(n576), .ZN(n511) );
  OAI221_X1 U65 ( .B1(n563), .B2(n29), .C1(n557), .C2(n22), .A(n577), .ZN(n518) );
  OAI221_X1 U66 ( .B1(n563), .B2(n12), .C1(n556), .C2(n5), .A(n576), .ZN(n501)
         );
  OAI221_X1 U67 ( .B1(n563), .B2(n19), .C1(n557), .C2(n12), .A(n576), .ZN(n508) );
  OAI221_X1 U68 ( .B1(n563), .B2(n54), .C1(n558), .C2(n47), .A(n577), .ZN(n543) );
  OAI221_X1 U69 ( .B1(n562), .B2(n9), .C1(n556), .C2(n2), .A(n576), .ZN(n498)
         );
  OAI221_X1 U70 ( .B1(n563), .B2(n16), .C1(n557), .C2(n9), .A(n576), .ZN(n505)
         );
  OAI221_X1 U71 ( .B1(n563), .B2(n13), .C1(n557), .C2(n6), .A(n576), .ZN(n502)
         );
  OAI221_X1 U72 ( .B1(n562), .B2(n20), .C1(n557), .C2(n13), .A(n576), .ZN(n509) );
  OAI221_X1 U73 ( .B1(n563), .B2(n48), .C1(n557), .C2(n41), .A(n577), .ZN(n537) );
  OAI221_X1 U74 ( .B1(n567), .B2(n31), .C1(n557), .C2(n24), .A(n577), .ZN(n520) );
  OAI221_X1 U75 ( .B1(n187), .B2(n53), .C1(n558), .C2(n46), .A(n577), .ZN(n542) );
  OAI221_X1 U76 ( .B1(n187), .B2(n50), .C1(n558), .C2(n43), .A(n577), .ZN(n539) );
  OAI221_X1 U77 ( .B1(n187), .B2(n26), .C1(n557), .C2(n19), .A(n577), .ZN(n515) );
  OAI221_X1 U78 ( .B1(n187), .B2(n51), .C1(n558), .C2(n44), .A(n577), .ZN(n540) );
  OAI221_X1 U79 ( .B1(n187), .B2(n27), .C1(n557), .C2(n20), .A(n577), .ZN(n516) );
  OAI221_X1 U80 ( .B1(n205), .B2(n565), .C1(n555), .C2(n103), .A(n575), .ZN(
        n476) );
  OAI221_X1 U81 ( .B1(n219), .B2(n562), .C1(n556), .C2(n117), .A(n575), .ZN(
        n490) );
  OAI221_X1 U82 ( .B1(n216), .B2(n563), .C1(n555), .C2(n114), .A(n575), .ZN(
        n487) );
  OAI221_X1 U83 ( .B1(n220), .B2(n565), .C1(n556), .C2(n118), .A(n575), .ZN(
        n491) );
  OAI221_X1 U84 ( .B1(n621), .B2(n564), .C1(n556), .C2(n121), .A(n575), .ZN(
        n494) );
  INV_X1 U85 ( .A(n223), .ZN(n621) );
  OAI221_X1 U86 ( .B1(n620), .B2(n566), .C1(n556), .C2(n120), .A(n575), .ZN(
        n493) );
  INV_X1 U87 ( .A(n222), .ZN(n620) );
  OAI22_X1 U88 ( .A1(n185), .A2(n141), .B1(n564), .B2(n154), .ZN(n390) );
  OAI22_X1 U89 ( .A1(n129), .A2(n142), .B1(n564), .B2(n155), .ZN(n391) );
  OAI22_X1 U90 ( .A1(n129), .A2(n144), .B1(n564), .B2(n157), .ZN(n393) );
  OAI22_X1 U91 ( .A1(n129), .A2(n38), .B1(n564), .B2(n45), .ZN(n534) );
  OAI22_X1 U92 ( .A1(n185), .A2(n35), .B1(n564), .B2(n42), .ZN(n531) );
  OAI22_X1 U93 ( .A1(n129), .A2(n11), .B1(n564), .B2(n18), .ZN(n507) );
  OAI22_X1 U94 ( .A1(n185), .A2(n39), .B1(n564), .B2(n46), .ZN(n535) );
  OAI22_X1 U95 ( .A1(n129), .A2(n36), .B1(n564), .B2(n43), .ZN(n532) );
  OAI22_X1 U96 ( .A1(n185), .A2(n40), .B1(n564), .B2(n47), .ZN(n536) );
  OAI22_X1 U97 ( .A1(n185), .A2(n37), .B1(n564), .B2(n44), .ZN(n533) );
  OAI22_X1 U98 ( .A1(n129), .A2(n34), .B1(n564), .B2(n41), .ZN(n530) );
  OAI22_X1 U99 ( .A1(n185), .A2(n48), .B1(n564), .B2(n55), .ZN(n544) );
  OAI22_X1 U100 ( .A1(n125), .A2(n165), .B1(n565), .B2(n178), .ZN(n414) );
  OAI22_X1 U101 ( .A1(n125), .A2(n166), .B1(n565), .B2(n179), .ZN(n415) );
  OAI22_X1 U102 ( .A1(n125), .A2(n167), .B1(n566), .B2(n180), .ZN(n416) );
  OAI22_X1 U103 ( .A1(n127), .A2(n161), .B1(n565), .B2(n174), .ZN(n410) );
  OAI22_X1 U104 ( .A1(n125), .A2(n168), .B1(n566), .B2(n181), .ZN(n417) );
  OAI22_X1 U105 ( .A1(n125), .A2(n169), .B1(n566), .B2(n182), .ZN(n418) );
  OAI22_X1 U106 ( .A1(n125), .A2(n170), .B1(n566), .B2(n183), .ZN(n419) );
  OAI22_X1 U107 ( .A1(n125), .A2(n164), .B1(n565), .B2(n177), .ZN(n413) );
  OAI22_X1 U108 ( .A1(n125), .A2(n171), .B1(n566), .B2(n184), .ZN(n420) );
  OAI22_X1 U109 ( .A1(n82), .A2(n60), .B1(n566), .B2(n89), .ZN(n438) );
  OAI22_X1 U110 ( .A1(n84), .A2(n74), .B1(n567), .B2(n103), .ZN(n452) );
  OAI22_X1 U111 ( .A1(n127), .A2(n59), .B1(n566), .B2(n88), .ZN(n437) );
  OAI22_X1 U112 ( .A1(n84), .A2(n73), .B1(n567), .B2(n102), .ZN(n451) );
  OAI22_X1 U113 ( .A1(n82), .A2(n58), .B1(n566), .B2(n87), .ZN(n436) );
  OAI22_X1 U114 ( .A1(n84), .A2(n72), .B1(n567), .B2(n101), .ZN(n450) );
  OAI22_X1 U115 ( .A1(n82), .A2(n62), .B1(n566), .B2(n91), .ZN(n440) );
  OAI22_X1 U116 ( .A1(n82), .A2(n71), .B1(n567), .B2(n100), .ZN(n449) );
  OAI22_X1 U117 ( .A1(n84), .A2(n75), .B1(n567), .B2(n104), .ZN(n453) );
  OAI22_X1 U118 ( .A1(n84), .A2(n83), .B1(n567), .B2(n108), .ZN(n457) );
  OAI22_X1 U119 ( .A1(n82), .A2(n69), .B1(n567), .B2(n98), .ZN(n447) );
  OAI22_X1 U120 ( .A1(n84), .A2(n81), .B1(n567), .B2(n107), .ZN(n456) );
  OAI22_X1 U121 ( .A1(n82), .A2(n68), .B1(n567), .B2(n97), .ZN(n446) );
  OAI22_X1 U122 ( .A1(n84), .A2(n79), .B1(n567), .B2(n106), .ZN(n455) );
  OAI22_X1 U123 ( .A1(n84), .A2(n77), .B1(n567), .B2(n105), .ZN(n454) );
  OAI22_X1 U124 ( .A1(n82), .A2(n66), .B1(n566), .B2(n95), .ZN(n444) );
  OAI22_X1 U125 ( .A1(n82), .A2(n56), .B1(n566), .B2(n85), .ZN(n434) );
  OAI22_X1 U126 ( .A1(n82), .A2(n70), .B1(n567), .B2(n99), .ZN(n448) );
  OAI22_X1 U127 ( .A1(n185), .A2(n31), .B1(n565), .B2(n38), .ZN(n527) );
  OAI22_X1 U128 ( .A1(n185), .A2(n21), .B1(n566), .B2(n28), .ZN(n517) );
  OAI22_X1 U129 ( .A1(n127), .A2(n28), .B1(n565), .B2(n35), .ZN(n524) );
  OAI22_X1 U130 ( .A1(n127), .A2(n18), .B1(n567), .B2(n25), .ZN(n514) );
  OAI22_X1 U131 ( .A1(n185), .A2(n25), .B1(n565), .B2(n32), .ZN(n521) );
  OAI22_X1 U132 ( .A1(n129), .A2(n32), .B1(n565), .B2(n39), .ZN(n528) );
  OAI22_X1 U133 ( .A1(n185), .A2(n29), .B1(n565), .B2(n36), .ZN(n525) );
  OAI22_X1 U134 ( .A1(n129), .A2(n26), .B1(n565), .B2(n33), .ZN(n522) );
  OAI22_X1 U135 ( .A1(n129), .A2(n33), .B1(n565), .B2(n40), .ZN(n529) );
  OAI22_X1 U136 ( .A1(n129), .A2(n23), .B1(n566), .B2(n30), .ZN(n519) );
  OAI22_X1 U137 ( .A1(n129), .A2(n30), .B1(n565), .B2(n37), .ZN(n526) );
  OAI22_X1 U138 ( .A1(n185), .A2(n27), .B1(n565), .B2(n34), .ZN(n523) );
  OAI221_X1 U139 ( .B1(n197), .B2(n562), .C1(n552), .C2(n180), .A(n572), .ZN(
        n429) );
  OAI221_X1 U140 ( .B1(n198), .B2(n564), .C1(n552), .C2(n181), .A(n572), .ZN(
        n430) );
  OAI221_X1 U141 ( .B1(n200), .B2(n563), .C1(n553), .C2(n183), .A(n572), .ZN(
        n432) );
  OAI221_X1 U142 ( .B1(n204), .B2(n564), .C1(n555), .C2(n102), .A(n574), .ZN(
        n475) );
  OAI221_X1 U143 ( .B1(n218), .B2(n565), .C1(n556), .C2(n116), .A(n575), .ZN(
        n489) );
  OAI221_X1 U144 ( .B1(n203), .B2(n566), .C1(n555), .C2(n101), .A(n574), .ZN(
        n474) );
  OAI221_X1 U145 ( .B1(n202), .B2(n567), .C1(n555), .C2(n100), .A(n574), .ZN(
        n473) );
  OAI221_X1 U146 ( .B1(n206), .B2(n559), .C1(n555), .C2(n104), .A(n575), .ZN(
        n477) );
  OAI221_X1 U147 ( .B1(n622), .B2(n560), .C1(n556), .C2(n122), .A(n575), .ZN(
        n495) );
  INV_X1 U148 ( .A(n224), .ZN(n622) );
  OAI221_X1 U149 ( .B1(n619), .B2(n561), .C1(n556), .C2(n119), .A(n575), .ZN(
        n492) );
  INV_X1 U150 ( .A(n221), .ZN(n619) );
  OAI221_X1 U151 ( .B1(n229), .B2(n563), .C1(n558), .C2(n52), .A(n578), .ZN(
        n548) );
  OAI221_X1 U152 ( .B1(n226), .B2(n562), .C1(n558), .C2(n49), .A(n577), .ZN(
        n545) );
  OAI221_X1 U153 ( .B1(n231), .B2(n564), .C1(n553), .C2(n54), .A(n578), .ZN(
        n550) );
  OAI221_X1 U154 ( .B1(n623), .B2(n564), .C1(n556), .C2(n123), .A(n575), .ZN(
        n496) );
  INV_X1 U155 ( .A(n225), .ZN(n623) );
  OAI221_X1 U156 ( .B1(n559), .B2(n152), .C1(n552), .C2(n139), .A(n570), .ZN(
        n388) );
  OAI221_X1 U157 ( .B1(n560), .B2(n165), .C1(n186), .C2(n152), .A(n571), .ZN(
        n401) );
  OAI221_X1 U158 ( .B1(n559), .B2(n146), .C1(n553), .C2(n133), .A(n570), .ZN(
        n382) );
  OAI221_X1 U159 ( .B1(n560), .B2(n159), .C1(n186), .C2(n146), .A(n571), .ZN(
        n395) );
  OAI221_X1 U160 ( .B1(n560), .B2(n172), .C1(n552), .C2(n159), .A(n572), .ZN(
        n408) );
  OAI221_X1 U161 ( .B1(n560), .B2(n153), .C1(n140), .C2(n82), .A(n571), .ZN(
        n389) );
  OAI221_X1 U162 ( .B1(n560), .B2(n166), .C1(n552), .C2(n153), .A(n571), .ZN(
        n402) );
  OAI221_X1 U163 ( .B1(n559), .B2(n147), .C1(n553), .C2(n134), .A(n570), .ZN(
        n383) );
  OAI221_X1 U164 ( .B1(n560), .B2(n160), .C1(n552), .C2(n147), .A(n571), .ZN(
        n396) );
  OAI221_X1 U165 ( .B1(n559), .B2(n173), .C1(n186), .C2(n160), .A(n572), .ZN(
        n409) );
  OAI221_X1 U166 ( .B1(n559), .B2(n141), .C1(n553), .C2(n126), .A(n570), .ZN(
        n377) );
  OAI221_X1 U167 ( .B1(n560), .B2(n167), .C1(n186), .C2(n154), .A(n571), .ZN(
        n403) );
  OAI221_X1 U168 ( .B1(n559), .B2(n148), .C1(n553), .C2(n135), .A(n570), .ZN(
        n384) );
  OAI221_X1 U169 ( .B1(n560), .B2(n161), .C1(n186), .C2(n148), .A(n571), .ZN(
        n397) );
  OAI221_X1 U170 ( .B1(n559), .B2(n142), .C1(n553), .C2(n128), .A(n570), .ZN(
        n378) );
  OAI221_X1 U171 ( .B1(n561), .B2(n168), .C1(n186), .C2(n155), .A(n572), .ZN(
        n404) );
  OAI221_X1 U172 ( .B1(n559), .B2(n149), .C1(n553), .C2(n136), .A(n570), .ZN(
        n385) );
  OAI221_X1 U173 ( .B1(n560), .B2(n162), .C1(n186), .C2(n149), .A(n571), .ZN(
        n398) );
  OAI221_X1 U174 ( .B1(n562), .B2(n175), .C1(n552), .C2(n162), .A(n572), .ZN(
        n411) );
  OAI221_X1 U175 ( .B1(n559), .B2(n143), .C1(n553), .C2(n130), .A(n570), .ZN(
        n379) );
  OAI221_X1 U176 ( .B1(n560), .B2(n156), .C1(n552), .C2(n143), .A(n571), .ZN(
        n392) );
  OAI221_X1 U177 ( .B1(n563), .B2(n169), .C1(n186), .C2(n156), .A(n572), .ZN(
        n405) );
  OAI221_X1 U178 ( .B1(n559), .B2(n150), .C1(n552), .C2(n137), .A(n570), .ZN(
        n386) );
  OAI221_X1 U179 ( .B1(n560), .B2(n163), .C1(n186), .C2(n150), .A(n571), .ZN(
        n399) );
  OAI221_X1 U180 ( .B1(n565), .B2(n176), .C1(n552), .C2(n163), .A(n572), .ZN(
        n412) );
  OAI221_X1 U181 ( .B1(n559), .B2(n144), .C1(n553), .C2(n131), .A(n570), .ZN(
        n380) );
  OAI221_X1 U182 ( .B1(n567), .B2(n170), .C1(n552), .C2(n157), .A(n572), .ZN(
        n406) );
  OAI221_X1 U183 ( .B1(n559), .B2(n151), .C1(n552), .C2(n138), .A(n570), .ZN(
        n387) );
  OAI221_X1 U184 ( .B1(n560), .B2(n164), .C1(n186), .C2(n151), .A(n571), .ZN(
        n400) );
  OAI221_X1 U185 ( .B1(n559), .B2(n145), .C1(n553), .C2(n132), .A(n570), .ZN(
        n381) );
  OAI221_X1 U186 ( .B1(n560), .B2(n158), .C1(n186), .C2(n145), .A(n571), .ZN(
        n394) );
  OAI221_X1 U187 ( .B1(n560), .B2(n171), .C1(n552), .C2(n158), .A(n572), .ZN(
        n407) );
  OAI221_X1 U188 ( .B1(n559), .B2(n93), .C1(n554), .C2(n64), .A(n573), .ZN(
        n442) );
  OAI221_X1 U189 ( .B1(n561), .B2(n92), .C1(n554), .C2(n63), .A(n573), .ZN(
        n441) );
  OAI221_X1 U190 ( .B1(n562), .B2(n86), .C1(n553), .C2(n57), .A(n572), .ZN(
        n435) );
  OAI221_X1 U191 ( .B1(n563), .B2(n90), .C1(n554), .C2(n61), .A(n573), .ZN(
        n439) );
  OAI22_X1 U192 ( .A1(n84), .A2(n178), .B1(n195), .B2(n559), .ZN(n427) );
  OAI22_X1 U193 ( .A1(n125), .A2(n172), .B1(n626), .B2(n560), .ZN(n421) );
  INV_X1 U194 ( .A(n189), .ZN(n626) );
  OAI22_X1 U195 ( .A1(n84), .A2(n179), .B1(n196), .B2(n561), .ZN(n428) );
  OAI22_X1 U196 ( .A1(n125), .A2(n173), .B1(n625), .B2(n562), .ZN(n422) );
  INV_X1 U197 ( .A(n190), .ZN(n625) );
  OAI22_X1 U198 ( .A1(n125), .A2(n175), .B1(n192), .B2(n563), .ZN(n424) );
  OAI22_X1 U199 ( .A1(n84), .A2(n182), .B1(n199), .B2(n565), .ZN(n431) );
  OAI22_X1 U200 ( .A1(n82), .A2(n184), .B1(n201), .B2(n187), .ZN(n433) );
  OAI22_X1 U201 ( .A1(n127), .A2(n113), .B1(n215), .B2(n187), .ZN(n486) );
  OAI22_X1 U202 ( .A1(n127), .A2(n112), .B1(n214), .B2(n187), .ZN(n485) );
  OAI22_X1 U203 ( .A1(n127), .A2(n111), .B1(n213), .B2(n187), .ZN(n484) );
  OAI22_X1 U204 ( .A1(n125), .A2(n105), .B1(n207), .B2(n187), .ZN(n478) );
  OAI22_X1 U205 ( .A1(n127), .A2(n109), .B1(n211), .B2(n187), .ZN(n482) );
  OAI22_X1 U206 ( .A1(n125), .A2(n174), .B1(n624), .B2(n566), .ZN(n423) );
  INV_X1 U207 ( .A(n191), .ZN(n624) );
  OAI22_X1 U208 ( .A1(n84), .A2(n176), .B1(n193), .B2(n567), .ZN(n425) );
  OAI22_X1 U209 ( .A1(n84), .A2(n177), .B1(n194), .B2(n559), .ZN(n426) );
  OAI22_X1 U210 ( .A1(n127), .A2(n110), .B1(n212), .B2(n560), .ZN(n483) );
  OAI22_X1 U211 ( .A1(n127), .A2(n115), .B1(n217), .B2(n561), .ZN(n488) );
  OAI22_X1 U212 ( .A1(n127), .A2(n108), .B1(n210), .B2(n562), .ZN(n481) );
  OAI22_X1 U213 ( .A1(n127), .A2(n107), .B1(n209), .B2(n563), .ZN(n480) );
  OAI22_X1 U214 ( .A1(n127), .A2(n106), .B1(n208), .B2(n564), .ZN(n479) );
  OAI22_X1 U215 ( .A1(n186), .A2(n53), .B1(n230), .B2(n567), .ZN(n549) );
  OAI22_X1 U216 ( .A1(n185), .A2(n50), .B1(n227), .B2(n566), .ZN(n546) );
  OAI22_X1 U217 ( .A1(n186), .A2(n51), .B1(n228), .B2(n559), .ZN(n547) );
  OAI22_X1 U218 ( .A1(n82), .A2(n55), .B1(n232), .B2(n560), .ZN(n551) );
  NAND2_X1 U219 ( .A1(ce), .A2(n578), .ZN(n187) );
  OAI22_X1 U220 ( .A1(n129), .A2(n14), .B1(n561), .B2(n21), .ZN(n510) );
  OAI22_X1 U221 ( .A1(n129), .A2(n16), .B1(n565), .B2(n23), .ZN(n512) );
  OAI22_X1 U222 ( .A1(n185), .A2(n17), .B1(n566), .B2(n24), .ZN(n513) );
  BUF_X1 U223 ( .A(rstn), .Z(n569) );
  NOR2_X1 U224 ( .A1(n610), .A2(n372), .ZN(N246) );
  XNOR2_X1 U225 ( .A(z1_next[63]), .B(n244), .ZN(n373) );
  XNOR2_X1 U226 ( .A(n164), .B(n375), .ZN(n374) );
  NOR2_X1 U227 ( .A1(n610), .A2(n368), .ZN(N247) );
  XNOR2_X1 U228 ( .A(z2_next[40]), .B(n225), .ZN(n369) );
  XNOR2_X1 U229 ( .A(n144), .B(n371), .ZN(n370) );
  NOR2_X1 U230 ( .A1(n609), .A2(n364), .ZN(N248) );
  XNOR2_X1 U231 ( .A(z2_next[41]), .B(n224), .ZN(n365) );
  XNOR2_X1 U232 ( .A(n143), .B(n367), .ZN(n366) );
  NOR2_X1 U233 ( .A1(n609), .A2(n360), .ZN(N249) );
  XNOR2_X1 U234 ( .A(n142), .B(n363), .ZN(n362) );
  XNOR2_X1 U235 ( .A(z2_next[42]), .B(n223), .ZN(n361) );
  NOR2_X1 U236 ( .A1(n608), .A2(n356), .ZN(N250) );
  XNOR2_X1 U237 ( .A(z2_next[43]), .B(n222), .ZN(n357) );
  XNOR2_X1 U238 ( .A(n141), .B(n359), .ZN(n358) );
  NOR2_X1 U239 ( .A1(n608), .A2(n352), .ZN(N251) );
  XNOR2_X1 U240 ( .A(z2_next[44]), .B(n221), .ZN(n353) );
  XNOR2_X1 U241 ( .A(n140), .B(n355), .ZN(n354) );
  NOR2_X1 U242 ( .A1(n607), .A2(n349), .ZN(N252) );
  XNOR2_X1 U243 ( .A(z3_next[37]), .B(z3_next[61]), .ZN(n350) );
  NOR2_X1 U244 ( .A1(n607), .A2(n346), .ZN(N253) );
  XNOR2_X1 U245 ( .A(z3_next[38]), .B(z3_next[62]), .ZN(n347) );
  NOR2_X1 U246 ( .A1(n606), .A2(n343), .ZN(N254) );
  XNOR2_X1 U247 ( .A(z3_next[39]), .B(z3_next[63]), .ZN(n344) );
  NOR2_X1 U248 ( .A1(n602), .A2(n327), .ZN(N262) );
  XNOR2_X1 U249 ( .A(n328), .B(n210), .ZN(n327) );
  XNOR2_X1 U250 ( .A(z3_next[16]), .B(n191), .ZN(n328) );
  NOR2_X1 U251 ( .A1(n602), .A2(n325), .ZN(N263) );
  XNOR2_X1 U252 ( .A(n326), .B(n209), .ZN(n325) );
  XNOR2_X1 U253 ( .A(z3_next[17]), .B(n190), .ZN(n326) );
  NOR2_X1 U254 ( .A1(n601), .A2(n323), .ZN(N264) );
  XNOR2_X1 U255 ( .A(n324), .B(n208), .ZN(n323) );
  XNOR2_X1 U256 ( .A(z3_next[18]), .B(n189), .ZN(n324) );
  NOR2_X1 U257 ( .A1(n601), .A2(n321), .ZN(N265) );
  XNOR2_X1 U258 ( .A(n322), .B(n207), .ZN(n321) );
  XNOR2_X1 U259 ( .A(z2_next[19]), .B(z3_next[19]), .ZN(n322) );
  NOR2_X1 U260 ( .A1(n600), .A2(n319), .ZN(N266) );
  XNOR2_X1 U261 ( .A(n320), .B(n206), .ZN(n319) );
  XNOR2_X1 U262 ( .A(z2_next[20]), .B(z3_next[20]), .ZN(n320) );
  NOR2_X1 U263 ( .A1(n600), .A2(n317), .ZN(N267) );
  XNOR2_X1 U264 ( .A(n318), .B(n205), .ZN(n317) );
  XNOR2_X1 U265 ( .A(z2_next[21]), .B(z3_next[21]), .ZN(n318) );
  NOR2_X1 U266 ( .A1(n599), .A2(n315), .ZN(N268) );
  XNOR2_X1 U267 ( .A(n316), .B(n204), .ZN(n315) );
  XNOR2_X1 U268 ( .A(z2_next[22]), .B(z3_next[22]), .ZN(n316) );
  NOR2_X1 U269 ( .A1(n599), .A2(n313), .ZN(N269) );
  XNOR2_X1 U270 ( .A(n314), .B(n203), .ZN(n313) );
  XNOR2_X1 U271 ( .A(z2_next[23]), .B(z3_next[23]), .ZN(n314) );
  NOR2_X1 U272 ( .A1(n598), .A2(n311), .ZN(N270) );
  XNOR2_X1 U273 ( .A(n312), .B(n202), .ZN(n311) );
  XNOR2_X1 U274 ( .A(z2_next[24]), .B(z3_next[24]), .ZN(n312) );
  NOR2_X1 U275 ( .A1(n598), .A2(n3090), .ZN(N271) );
  XNOR2_X1 U276 ( .A(z1_next[25]), .B(n310), .ZN(n3090) );
  XNOR2_X1 U277 ( .A(n46), .B(z2_next[25]), .ZN(n310) );
  NOR2_X1 U278 ( .A1(n597), .A2(n3070), .ZN(N272) );
  XNOR2_X1 U279 ( .A(z1_next[26]), .B(n3080), .ZN(n3070) );
  XNOR2_X1 U280 ( .A(n45), .B(z2_next[26]), .ZN(n3080) );
  NOR2_X1 U281 ( .A1(n597), .A2(n3050), .ZN(N273) );
  XNOR2_X1 U282 ( .A(z1_next[27]), .B(n3060), .ZN(n3050) );
  XNOR2_X1 U283 ( .A(n44), .B(z2_next[27]), .ZN(n3060) );
  NOR2_X1 U284 ( .A1(n596), .A2(n3030), .ZN(N274) );
  XNOR2_X1 U285 ( .A(z1_next[28]), .B(n3040), .ZN(n3030) );
  XNOR2_X1 U286 ( .A(n43), .B(z2_next[28]), .ZN(n3040) );
  NOR2_X1 U287 ( .A1(n596), .A2(n3010), .ZN(N275) );
  XNOR2_X1 U288 ( .A(z1_next[29]), .B(n3020), .ZN(n3010) );
  XNOR2_X1 U289 ( .A(n42), .B(z2_next[29]), .ZN(n3020) );
  NOR2_X1 U290 ( .A1(n595), .A2(n2990), .ZN(N276) );
  XNOR2_X1 U291 ( .A(z1_next[30]), .B(n3000), .ZN(n2990) );
  XNOR2_X1 U292 ( .A(n41), .B(z2_next[30]), .ZN(n3000) );
  NOR2_X1 U293 ( .A1(n595), .A2(n2970), .ZN(N277) );
  XNOR2_X1 U294 ( .A(z1_next[31]), .B(n2980), .ZN(n2970) );
  XNOR2_X1 U295 ( .A(n40), .B(z2_next[31]), .ZN(n2980) );
  NOR2_X1 U296 ( .A1(n594), .A2(n2950), .ZN(N278) );
  XNOR2_X1 U297 ( .A(z1_next[32]), .B(n2960), .ZN(n2950) );
  XNOR2_X1 U298 ( .A(n39), .B(z2_next[32]), .ZN(n2960) );
  NOR2_X1 U299 ( .A1(n594), .A2(n2930), .ZN(N279) );
  XNOR2_X1 U300 ( .A(z1_next[33]), .B(n2940), .ZN(n2930) );
  XNOR2_X1 U301 ( .A(n38), .B(z2_next[33]), .ZN(n2940) );
  NOR2_X1 U302 ( .A1(n593), .A2(n2910), .ZN(N280) );
  XNOR2_X1 U303 ( .A(z1_next[34]), .B(n2920), .ZN(n2910) );
  XNOR2_X1 U304 ( .A(n37), .B(z2_next[34]), .ZN(n2920) );
  NOR2_X1 U305 ( .A1(n593), .A2(n2890), .ZN(N281) );
  XNOR2_X1 U306 ( .A(z1_next[35]), .B(n2900), .ZN(n2890) );
  XNOR2_X1 U307 ( .A(n36), .B(z2_next[35]), .ZN(n2900) );
  NOR2_X1 U308 ( .A1(n592), .A2(n2870), .ZN(N282) );
  XNOR2_X1 U309 ( .A(z1_next[36]), .B(n2880), .ZN(n2870) );
  XNOR2_X1 U310 ( .A(n35), .B(z2_next[36]), .ZN(n2880) );
  NOR2_X1 U311 ( .A1(n592), .A2(n2850), .ZN(N283) );
  XNOR2_X1 U312 ( .A(z1_next[37]), .B(n2860), .ZN(n2850) );
  XNOR2_X1 U313 ( .A(n34), .B(z2_next[37]), .ZN(n2860) );
  NOR2_X1 U314 ( .A1(n591), .A2(n2830), .ZN(N284) );
  XNOR2_X1 U315 ( .A(z1_next[38]), .B(n2840), .ZN(n2830) );
  XNOR2_X1 U316 ( .A(n33), .B(z2_next[38]), .ZN(n2840) );
  NOR2_X1 U317 ( .A1(n591), .A2(n2810), .ZN(N285) );
  XNOR2_X1 U318 ( .A(z1_next[39]), .B(n2820), .ZN(n2810) );
  XNOR2_X1 U319 ( .A(n32), .B(z2_next[39]), .ZN(n2820) );
  NOR2_X1 U320 ( .A1(n590), .A2(n2790), .ZN(N286) );
  XNOR2_X1 U321 ( .A(z1_next[40]), .B(n2800), .ZN(n2790) );
  XNOR2_X1 U322 ( .A(n31), .B(z2_next[40]), .ZN(n2800) );
  NOR2_X1 U323 ( .A1(n590), .A2(n2770), .ZN(N287) );
  XNOR2_X1 U324 ( .A(z1_next[41]), .B(n2780), .ZN(n2770) );
  XNOR2_X1 U325 ( .A(n30), .B(z2_next[41]), .ZN(n2780) );
  NOR2_X1 U326 ( .A1(n589), .A2(n2750), .ZN(N288) );
  XNOR2_X1 U327 ( .A(z1_next[42]), .B(n2760), .ZN(n2750) );
  XNOR2_X1 U328 ( .A(n29), .B(z2_next[42]), .ZN(n2760) );
  NOR2_X1 U329 ( .A1(n589), .A2(n2730), .ZN(N289) );
  XNOR2_X1 U330 ( .A(z1_next[43]), .B(n2740), .ZN(n2730) );
  XNOR2_X1 U331 ( .A(n28), .B(z2_next[43]), .ZN(n2740) );
  NOR2_X1 U332 ( .A1(n588), .A2(n2710), .ZN(N290) );
  XNOR2_X1 U333 ( .A(z1_next[44]), .B(n2720), .ZN(n2710) );
  XNOR2_X1 U334 ( .A(n27), .B(z2_next[44]), .ZN(n2720) );
  NOR2_X1 U335 ( .A1(n588), .A2(n2690), .ZN(N291) );
  XNOR2_X1 U336 ( .A(z1_next[45]), .B(n2700), .ZN(n2690) );
  XNOR2_X1 U337 ( .A(n26), .B(z2_next[45]), .ZN(n2700) );
  NOR2_X1 U338 ( .A1(n587), .A2(n2670), .ZN(N292) );
  XNOR2_X1 U339 ( .A(z1_next[46]), .B(n2680), .ZN(n2670) );
  XNOR2_X1 U340 ( .A(n25), .B(z2_next[46]), .ZN(n2680) );
  NOR2_X1 U341 ( .A1(n587), .A2(n2650), .ZN(N293) );
  XNOR2_X1 U342 ( .A(z1_next[47]), .B(n2660), .ZN(n2650) );
  XNOR2_X1 U343 ( .A(n24), .B(z2_next[47]), .ZN(n2660) );
  NOR2_X1 U344 ( .A1(n586), .A2(n2630), .ZN(N294) );
  XNOR2_X1 U345 ( .A(z1_next[48]), .B(n2640), .ZN(n2630) );
  XNOR2_X1 U346 ( .A(n23), .B(z2_next[48]), .ZN(n2640) );
  NOR2_X1 U347 ( .A1(n586), .A2(n2610), .ZN(N295) );
  XNOR2_X1 U348 ( .A(z1_next[49]), .B(n2620), .ZN(n2610) );
  XNOR2_X1 U349 ( .A(n22), .B(z2_next[49]), .ZN(n2620) );
  NOR2_X1 U350 ( .A1(n585), .A2(n2590), .ZN(N296) );
  XNOR2_X1 U351 ( .A(z1_next[50]), .B(n2600), .ZN(n2590) );
  XNOR2_X1 U352 ( .A(n21), .B(z2_next[50]), .ZN(n2600) );
  NOR2_X1 U353 ( .A1(n585), .A2(n2570), .ZN(N297) );
  XNOR2_X1 U354 ( .A(z1_next[51]), .B(n2580), .ZN(n2570) );
  XNOR2_X1 U355 ( .A(n20), .B(z2_next[51]), .ZN(n2580) );
  NOR2_X1 U356 ( .A1(n584), .A2(n2550), .ZN(N298) );
  XNOR2_X1 U357 ( .A(z1_next[52]), .B(n2560), .ZN(n2550) );
  XNOR2_X1 U358 ( .A(n19), .B(z2_next[52]), .ZN(n2560) );
  NOR2_X1 U359 ( .A1(n584), .A2(n2530), .ZN(N299) );
  XNOR2_X1 U360 ( .A(z1_next[53]), .B(n2540), .ZN(n2530) );
  XNOR2_X1 U361 ( .A(n18), .B(z2_next[53]), .ZN(n2540) );
  NOR2_X1 U362 ( .A1(n583), .A2(n2510), .ZN(N300) );
  XNOR2_X1 U363 ( .A(z1_next[54]), .B(n2520), .ZN(n2510) );
  XNOR2_X1 U364 ( .A(n17), .B(z2_next[54]), .ZN(n2520) );
  NOR2_X1 U365 ( .A1(n583), .A2(n2490), .ZN(N301) );
  XNOR2_X1 U366 ( .A(z1_next[55]), .B(n2500), .ZN(n2490) );
  XNOR2_X1 U367 ( .A(n16), .B(z2_next[55]), .ZN(n2500) );
  NOR2_X1 U368 ( .A1(n582), .A2(n2470), .ZN(N302) );
  XNOR2_X1 U369 ( .A(z1_next[56]), .B(n2480), .ZN(n2470) );
  XNOR2_X1 U370 ( .A(n15), .B(z2_next[56]), .ZN(n2480) );
  NOR2_X1 U371 ( .A1(n582), .A2(n245), .ZN(N303) );
  XNOR2_X1 U372 ( .A(z1_next[57]), .B(n2460), .ZN(n245) );
  XNOR2_X1 U373 ( .A(n14), .B(z2_next[57]), .ZN(n2460) );
  NOR2_X1 U374 ( .A1(n581), .A2(n243), .ZN(N304) );
  XNOR2_X1 U375 ( .A(z3_next[58]), .B(n244), .ZN(n243) );
  NOR2_X1 U376 ( .A1(n581), .A2(n241), .ZN(N305) );
  XNOR2_X1 U377 ( .A(z1_next[59]), .B(n242), .ZN(n241) );
  XNOR2_X1 U378 ( .A(n12), .B(z2_next[59]), .ZN(n242) );
  NOR2_X1 U379 ( .A1(n580), .A2(n239), .ZN(N306) );
  XNOR2_X1 U380 ( .A(z1_next[60]), .B(n240), .ZN(n239) );
  XNOR2_X1 U381 ( .A(n11), .B(z2_next[60]), .ZN(n240) );
  NOR2_X1 U382 ( .A1(n580), .A2(n237), .ZN(N307) );
  XNOR2_X1 U383 ( .A(z1_next[61]), .B(n238), .ZN(n237) );
  XNOR2_X1 U384 ( .A(n10), .B(z2_next[61]), .ZN(n238) );
  NOR2_X1 U385 ( .A1(n579), .A2(n235), .ZN(N308) );
  XNOR2_X1 U386 ( .A(z1_next[62]), .B(n236), .ZN(n235) );
  XNOR2_X1 U387 ( .A(n9), .B(z2_next[62]), .ZN(n236) );
  NOR2_X1 U388 ( .A1(n579), .A2(n233), .ZN(N309) );
  XNOR2_X1 U389 ( .A(z1_next[63]), .B(n234), .ZN(n233) );
  XNOR2_X1 U390 ( .A(n8), .B(z2_next[63]), .ZN(n234) );
  XNOR2_X1 U391 ( .A(n90), .B(z2_next[58]), .ZN(n244) );
  XNOR2_X1 U392 ( .A(n62), .B(n57), .ZN(n203) );
  XNOR2_X1 U393 ( .A(n64), .B(n59), .ZN(n205) );
  XNOR2_X1 U394 ( .A(n63), .B(n58), .ZN(n204) );
  XNOR2_X1 U395 ( .A(n61), .B(n56), .ZN(n202) );
  XNOR2_X1 U396 ( .A(n65), .B(n60), .ZN(n206) );
  XNOR2_X1 U397 ( .A(z1[40]), .B(n89), .ZN(n225) );
  XNOR2_X1 U398 ( .A(z1[41]), .B(n88), .ZN(n224) );
  XNOR2_X1 U399 ( .A(z1[42]), .B(n87), .ZN(n223) );
  XNOR2_X1 U400 ( .A(z1[44]), .B(n85), .ZN(n221) );
  XNOR2_X1 U401 ( .A(z1[43]), .B(n86), .ZN(n222) );
  XNOR2_X1 U402 ( .A(z2[61]), .B(n148), .ZN(n191) );
  XNOR2_X1 U403 ( .A(z2[62]), .B(n147), .ZN(n190) );
  XNOR2_X1 U404 ( .A(z2[63]), .B(n146), .ZN(n189) );
  XNOR2_X1 U405 ( .A(n67), .B(n62), .ZN(n208) );
  XNOR2_X1 U442 ( .A(n69), .B(n64), .ZN(n210) );
  XNOR2_X1 U443 ( .A(n68), .B(n63), .ZN(n209) );
  XNOR2_X1 U444 ( .A(n66), .B(n61), .ZN(n207) );
  XNOR2_X1 U445 ( .A(n138), .B(n157), .ZN(n200) );
  XNOR2_X1 U446 ( .A(n136), .B(n155), .ZN(n198) );
  XNOR2_X1 U447 ( .A(n135), .B(n154), .ZN(n197) );
  XNOR2_X1 U448 ( .A(z3[58]), .B(z3_next[41]), .ZN(n231) );
  XNOR2_X1 U449 ( .A(z3[60]), .B(z3_next[43]), .ZN(n229) );
  XNOR2_X1 U450 ( .A(z3[63]), .B(z3_next[46]), .ZN(n226) );
  XNOR2_X1 U451 ( .A(n139), .B(n158), .ZN(n201) );
  XNOR2_X1 U452 ( .A(n137), .B(n156), .ZN(n199) );
  XNOR2_X1 U453 ( .A(n134), .B(n153), .ZN(n196) );
  XNOR2_X1 U454 ( .A(n133), .B(n152), .ZN(n195) );
  XNOR2_X1 U455 ( .A(n132), .B(n151), .ZN(n194) );
  XNOR2_X1 U456 ( .A(n131), .B(n150), .ZN(n193) );
  XNOR2_X1 U457 ( .A(n130), .B(n149), .ZN(n192) );
  XNOR2_X1 U458 ( .A(z3[57]), .B(z3_next[40]), .ZN(n232) );
  XNOR2_X1 U459 ( .A(z3[59]), .B(z3_next[42]), .ZN(n230) );
  XNOR2_X1 U460 ( .A(z3[61]), .B(z3_next[44]), .ZN(n228) );
  XNOR2_X1 U461 ( .A(z3[62]), .B(z3_next[45]), .ZN(n227) );
  XNOR2_X1 U462 ( .A(n16), .B(z3_next[31]), .ZN(n375) );
  XNOR2_X1 U463 ( .A(n14), .B(z3_next[33]), .ZN(n367) );
  XNOR2_X1 U464 ( .A(n11), .B(z3_next[36]), .ZN(n355) );
  XNOR2_X1 U465 ( .A(n15), .B(z3_next[32]), .ZN(n371) );
  XNOR2_X1 U466 ( .A(n12), .B(z3_next[35]), .ZN(n359) );
  XNOR2_X1 U467 ( .A(n13), .B(z3_next[34]), .ZN(n363) );
  BUF_X1 U468 ( .A(n80), .Z(n558) );
  INV_X1 U469 ( .A(n568), .ZN(n561) );
  INV_X1 U470 ( .A(n568), .ZN(n562) );
  INV_X1 U471 ( .A(n568), .ZN(n563) );
  INV_X1 U472 ( .A(n568), .ZN(n564) );
  INV_X1 U473 ( .A(n568), .ZN(n565) );
  INV_X1 U474 ( .A(n568), .ZN(n566) );
  INV_X1 U475 ( .A(n568), .ZN(n567) );
  INV_X1 U476 ( .A(n613), .ZN(n578) );
  BUF_X1 U477 ( .A(n615), .Z(n579) );
  BUF_X1 U478 ( .A(n614), .Z(n580) );
  BUF_X1 U479 ( .A(n616), .Z(n581) );
  BUF_X1 U480 ( .A(n615), .Z(n582) );
  BUF_X1 U481 ( .A(n614), .Z(n583) );
  BUF_X1 U482 ( .A(n614), .Z(n584) );
  BUF_X1 U483 ( .A(n616), .Z(n585) );
  BUF_X1 U484 ( .A(n615), .Z(n586) );
  BUF_X1 U485 ( .A(n616), .Z(n587) );
  BUF_X1 U486 ( .A(n615), .Z(n588) );
  BUF_X1 U487 ( .A(n614), .Z(n589) );
  BUF_X1 U488 ( .A(n616), .Z(n590) );
  BUF_X1 U489 ( .A(n618), .Z(n591) );
  BUF_X1 U490 ( .A(n617), .Z(n592) );
  BUF_X1 U491 ( .A(n616), .Z(n593) );
  BUF_X1 U492 ( .A(n615), .Z(n594) );
  BUF_X1 U493 ( .A(n614), .Z(n595) );
  BUF_X1 U494 ( .A(n618), .Z(n596) );
  BUF_X1 U495 ( .A(n618), .Z(n597) );
  BUF_X1 U496 ( .A(n618), .Z(n598) );
  BUF_X1 U497 ( .A(n617), .Z(n599) );
  BUF_X1 U498 ( .A(n617), .Z(n600) );
  BUF_X1 U499 ( .A(n617), .Z(n601) );
  BUF_X1 U500 ( .A(n616), .Z(n602) );
  BUF_X1 U501 ( .A(n616), .Z(n603) );
  BUF_X1 U502 ( .A(n616), .Z(n604) );
  BUF_X1 U503 ( .A(n615), .Z(n605) );
  BUF_X1 U504 ( .A(n615), .Z(n606) );
  BUF_X1 U505 ( .A(n615), .Z(n607) );
  BUF_X1 U506 ( .A(n614), .Z(n608) );
  BUF_X1 U507 ( .A(n614), .Z(n609) );
  BUF_X1 U508 ( .A(n614), .Z(n610) );
  BUF_X1 U509 ( .A(n618), .Z(n611) );
  BUF_X1 U510 ( .A(n617), .Z(n612) );
  BUF_X1 U511 ( .A(n618), .Z(n613) );
  INV_X1 U512 ( .A(n569), .ZN(n614) );
  INV_X1 U513 ( .A(n569), .ZN(n615) );
  INV_X1 U514 ( .A(n569), .ZN(n616) );
  INV_X1 U515 ( .A(n569), .ZN(n617) );
  INV_X1 U516 ( .A(n569), .ZN(n618) );
endmodule


module gng_lzd ( data_in, data_out );
  input [60:0] data_in;
  output [5:0] data_out;
  wire   n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n1, n2, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41;

  NOR4_X2 U44 ( .A1(data_in[45]), .A2(n4), .A3(data_in[47]), .A4(data_in[46]), 
        .ZN(n55) );
  NOR4_X2 U76 ( .A1(data_in[13]), .A2(n23), .A3(data_in[15]), .A4(data_in[14]), 
        .ZN(n48) );
  NOR4_X1 U2 ( .A1(data_in[55]), .A2(data_in[56]), .A3(data_in[54]), .A4(n98), 
        .ZN(n45) );
  OAI222_X1 U3 ( .A1(n82), .A2(n47), .B1(n55), .B2(n83), .C1(n84), .C2(n42), 
        .ZN(data_out[0]) );
  NOR4_X1 U4 ( .A1(n85), .A2(n86), .A3(n87), .A4(n88), .ZN(n84) );
  NOR4_X1 U5 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(n83) );
  OAI221_X1 U6 ( .B1(data_out[5]), .B2(n59), .C1(n60), .C2(n43), .A(n61), .ZN(
        data_out[1]) );
  AOI222_X1 U7 ( .A1(n67), .A2(n37), .B1(n68), .B2(n35), .C1(n69), .C2(n40), 
        .ZN(n60) );
  AOI22_X1 U8 ( .A1(n55), .A2(n70), .B1(n71), .B2(n2), .ZN(n59) );
  OAI221_X1 U9 ( .B1(n33), .B2(n43), .C1(n14), .C2(n42), .A(n44), .ZN(
        data_out[3]) );
  AOI21_X1 U10 ( .B1(n45), .B2(n2), .A(n46), .ZN(n44) );
  NOR3_X1 U11 ( .A1(n47), .A2(n48), .A3(n24), .ZN(n46) );
  OAI22_X1 U12 ( .A1(data_out[5]), .A2(n49), .B1(n50), .B2(n47), .ZN(
        data_out[2]) );
  AOI22_X1 U13 ( .A1(n48), .A2(n51), .B1(n52), .B2(n22), .ZN(n50) );
  AOI22_X1 U14 ( .A1(n55), .A2(n56), .B1(n57), .B2(n2), .ZN(n49) );
  NAND2_X1 U15 ( .A1(n42), .A2(n43), .ZN(data_out[4]) );
  NAND2_X1 U16 ( .A1(n55), .A2(n47), .ZN(n42) );
  INV_X1 U17 ( .A(n55), .ZN(n2) );
  NAND2_X1 U18 ( .A1(data_out[5]), .A2(n48), .ZN(n43) );
  INV_X1 U19 ( .A(n48), .ZN(n22) );
  INV_X1 U20 ( .A(n45), .ZN(n5) );
  OAI22_X1 U21 ( .A1(n54), .A2(n34), .B1(n33), .B2(n39), .ZN(n51) );
  OAI22_X1 U22 ( .A1(n58), .A2(n15), .B1(n18), .B2(n14), .ZN(n56) );
  INV_X1 U23 ( .A(n53), .ZN(n24) );
  INV_X1 U24 ( .A(n54), .ZN(n33) );
  INV_X1 U25 ( .A(n58), .ZN(n14) );
  OAI22_X1 U26 ( .A1(n45), .A2(n6), .B1(n9), .B2(n5), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n53), .A2(n25), .B1(n30), .B2(n24), .ZN(n52) );
  INV_X1 U28 ( .A(n47), .ZN(data_out[5]) );
  INV_X1 U29 ( .A(n114), .ZN(n34) );
  INV_X1 U30 ( .A(n108), .ZN(n25) );
  INV_X1 U31 ( .A(n89), .ZN(n15) );
  INV_X1 U32 ( .A(n95), .ZN(n6) );
  INV_X1 U33 ( .A(n107), .ZN(n30) );
  INV_X1 U34 ( .A(n96), .ZN(n9) );
  INV_X1 U35 ( .A(n90), .ZN(n18) );
  INV_X1 U36 ( .A(n106), .ZN(n23) );
  INV_X1 U37 ( .A(n75), .ZN(n4) );
  INV_X1 U38 ( .A(n113), .ZN(n39) );
  OR2_X1 U39 ( .A1(data_in[53]), .A2(n6), .ZN(n98) );
  NOR4_X1 U40 ( .A1(data_in[7]), .A2(data_in[8]), .A3(data_in[6]), .A4(n115), 
        .ZN(n54) );
  OR2_X1 U41 ( .A1(data_in[5]), .A2(n34), .ZN(n115) );
  NOR4_X1 U42 ( .A1(data_in[23]), .A2(data_in[24]), .A3(data_in[22]), .A4(n116), .ZN(n53) );
  OR2_X1 U43 ( .A1(data_in[21]), .A2(n25), .ZN(n116) );
  NOR4_X1 U45 ( .A1(data_in[18]), .A2(data_in[17]), .A3(data_in[20]), .A4(
        data_in[19]), .ZN(n107) );
  NOR4_X1 U46 ( .A1(data_in[50]), .A2(data_in[49]), .A3(data_in[52]), .A4(
        data_in[51]), .ZN(n96) );
  NOR4_X1 U47 ( .A1(data_in[34]), .A2(data_in[33]), .A3(data_in[36]), .A4(
        data_in[35]), .ZN(n90) );
  NOR4_X1 U48 ( .A1(data_in[11]), .A2(data_in[10]), .A3(data_in[9]), .A4(
        data_in[12]), .ZN(n114) );
  NOR4_X1 U49 ( .A1(data_in[26]), .A2(data_in[25]), .A3(data_in[28]), .A4(
        data_in[27]), .ZN(n108) );
  NAND3_X1 U50 ( .A1(n80), .A2(n55), .A3(n97), .ZN(n47) );
  NOR3_X1 U51 ( .A1(data_in[29]), .A2(data_in[31]), .A3(data_in[30]), .ZN(n97)
         );
  NOR3_X1 U52 ( .A1(data_in[32]), .A2(n18), .A3(n14), .ZN(n80) );
  NOR4_X1 U53 ( .A1(data_in[42]), .A2(data_in[41]), .A3(data_in[44]), .A4(
        data_in[43]), .ZN(n89) );
  NOR4_X1 U54 ( .A1(data_in[58]), .A2(data_in[57]), .A3(data_in[60]), .A4(
        data_in[59]), .ZN(n95) );
  NOR3_X1 U55 ( .A1(data_in[48]), .A2(n9), .A3(n5), .ZN(n75) );
  NOR3_X1 U56 ( .A1(data_in[16]), .A2(n30), .A3(n24), .ZN(n106) );
  NOR3_X1 U57 ( .A1(n107), .A2(data_in[20]), .A3(n24), .ZN(n66) );
  NOR3_X1 U58 ( .A1(n53), .A2(data_in[24]), .A3(n25), .ZN(n63) );
  NOR3_X1 U59 ( .A1(n54), .A2(data_in[8]), .A3(n34), .ZN(n67) );
  NOR3_X1 U60 ( .A1(n96), .A2(data_in[52]), .A3(n5), .ZN(n76) );
  NOR3_X1 U61 ( .A1(n90), .A2(data_in[36]), .A3(n14), .ZN(n81) );
  NOR3_X1 U62 ( .A1(n113), .A2(data_in[4]), .A3(n33), .ZN(n69) );
  AOI22_X1 U63 ( .A1(n48), .A2(n100), .B1(n101), .B2(n22), .ZN(n82) );
  NAND4_X1 U64 ( .A1(n109), .A2(n110), .A3(n111), .A4(n112), .ZN(n100) );
  NAND4_X1 U65 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(n101) );
  OAI21_X1 U66 ( .B1(data_in[11]), .B2(n36), .A(n68), .ZN(n111) );
  OAI221_X1 U67 ( .B1(data_in[39]), .B2(n77), .C1(data_in[43]), .C2(n78), .A(
        n79), .ZN(n70) );
  AOI22_X1 U68 ( .A1(n80), .A2(n20), .B1(n81), .B2(n19), .ZN(n79) );
  OAI221_X1 U69 ( .B1(data_in[55]), .B2(n72), .C1(data_in[59]), .C2(n73), .A(
        n74), .ZN(n71) );
  AOI22_X1 U70 ( .A1(n75), .A2(n11), .B1(n76), .B2(n10), .ZN(n74) );
  OAI22_X1 U71 ( .A1(n23), .A2(data_in[15]), .B1(n21), .B2(data_in[19]), .ZN(
        n65) );
  INV_X1 U72 ( .A(n66), .ZN(n21) );
  AOI21_X1 U73 ( .B1(data_in[54]), .B2(n8), .A(n72), .ZN(n93) );
  INV_X1 U74 ( .A(data_in[55]), .ZN(n8) );
  AOI21_X1 U75 ( .B1(data_in[38]), .B2(n17), .A(n77), .ZN(n87) );
  INV_X1 U77 ( .A(data_in[39]), .ZN(n17) );
  AOI21_X1 U78 ( .B1(data_in[50]), .B2(n10), .A(n1), .ZN(n92) );
  INV_X1 U79 ( .A(n76), .ZN(n1) );
  AOI21_X1 U80 ( .B1(data_in[34]), .B2(n19), .A(n12), .ZN(n86) );
  INV_X1 U81 ( .A(n81), .ZN(n12) );
  AOI21_X1 U82 ( .B1(data_in[46]), .B2(n11), .A(n4), .ZN(n91) );
  AOI21_X1 U83 ( .B1(data_in[30]), .B2(n20), .A(n13), .ZN(n85) );
  INV_X1 U84 ( .A(n80), .ZN(n13) );
  OAI21_X1 U85 ( .B1(data_in[15]), .B2(n32), .A(n106), .ZN(n105) );
  INV_X1 U86 ( .A(data_in[14]), .ZN(n32) );
  OAI21_X1 U87 ( .B1(data_in[19]), .B2(n31), .A(n66), .ZN(n104) );
  INV_X1 U88 ( .A(data_in[18]), .ZN(n31) );
  OAI21_X1 U89 ( .B1(data_in[3]), .B2(n41), .A(n69), .ZN(n110) );
  INV_X1 U90 ( .A(data_in[2]), .ZN(n41) );
  OAI21_X1 U91 ( .B1(data_in[23]), .B2(n29), .A(n63), .ZN(n103) );
  INV_X1 U92 ( .A(data_in[22]), .ZN(n29) );
  OAI21_X1 U93 ( .B1(data_in[7]), .B2(n38), .A(n67), .ZN(n109) );
  INV_X1 U94 ( .A(data_in[6]), .ZN(n38) );
  OR3_X1 U95 ( .A1(n45), .A2(data_in[56]), .A3(n6), .ZN(n72) );
  OR3_X1 U96 ( .A1(n58), .A2(data_in[40]), .A3(n15), .ZN(n77) );
  OR3_X1 U97 ( .A1(data_in[0]), .A2(n33), .A3(n39), .ZN(n112) );
  OR3_X1 U98 ( .A1(n62), .A2(n48), .A3(n47), .ZN(n61) );
  AOI221_X1 U99 ( .B1(n28), .B2(n63), .C1(n26), .C2(n64), .A(n65), .ZN(n62) );
  INV_X1 U100 ( .A(data_in[27]), .ZN(n26) );
  INV_X1 U101 ( .A(data_in[23]), .ZN(n28) );
  NOR4_X1 U102 ( .A1(data_in[39]), .A2(data_in[40]), .A3(data_in[38]), .A4(n99), .ZN(n58) );
  OR2_X1 U103 ( .A1(data_in[37]), .A2(n15), .ZN(n99) );
  NOR4_X1 U104 ( .A1(data_in[2]), .A2(data_in[1]), .A3(data_in[4]), .A4(
        data_in[3]), .ZN(n113) );
  NOR2_X1 U105 ( .A1(n108), .A2(data_in[28]), .ZN(n64) );
  NOR2_X1 U106 ( .A1(n114), .A2(data_in[12]), .ZN(n68) );
  AOI21_X1 U107 ( .B1(data_in[58]), .B2(n7), .A(n73), .ZN(n94) );
  INV_X1 U108 ( .A(data_in[59]), .ZN(n7) );
  AOI21_X1 U109 ( .B1(data_in[42]), .B2(n16), .A(n78), .ZN(n88) );
  INV_X1 U110 ( .A(data_in[43]), .ZN(n16) );
  OAI21_X1 U111 ( .B1(data_in[27]), .B2(n27), .A(n64), .ZN(n102) );
  INV_X1 U112 ( .A(data_in[26]), .ZN(n27) );
  OR2_X1 U113 ( .A1(n95), .A2(data_in[60]), .ZN(n73) );
  OR2_X1 U114 ( .A1(n89), .A2(data_in[44]), .ZN(n78) );
  INV_X1 U115 ( .A(data_in[51]), .ZN(n10) );
  INV_X1 U116 ( .A(data_in[35]), .ZN(n19) );
  INV_X1 U117 ( .A(data_in[47]), .ZN(n11) );
  INV_X1 U118 ( .A(data_in[31]), .ZN(n20) );
  INV_X1 U119 ( .A(data_in[3]), .ZN(n40) );
  INV_X1 U120 ( .A(data_in[11]), .ZN(n35) );
  INV_X1 U121 ( .A(data_in[7]), .ZN(n37) );
  INV_X1 U122 ( .A(data_in[10]), .ZN(n36) );
endmodule


module gng_coef ( clk, addr, c0, c1, c2 );
  input [7:0] addr;
  output [17:0] c0;
  output [17:0] c1;
  output [16:0] c2;
  input clk;
  wire   N464, N468, N487, N509, N1318, N1333, N1352, N1952, N1975, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n13180,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n13330, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n13520, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n408, n409, n410, n411, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n4640, n465, n466, n467, n4680, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n4870, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n5090, n510, n511, n512, n513, n514, n515, n516, n1499,
         n1500, n1501, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
  wire   [48:0] d;

  DFF_X1 c2_reg_16_ ( .D(N1952), .CK(clk), .Q(c2[16]) );
  DFF_X1 c2_reg_15_ ( .D(N1975), .CK(clk), .Q(c2[15]) );
  DFF_X1 c2_reg_14_ ( .D(d[14]), .CK(clk), .Q(c2[14]) );
  DFF_X1 c2_reg_13_ ( .D(d[13]), .CK(clk), .Q(c2[13]) );
  DFF_X1 c2_reg_12_ ( .D(d[12]), .CK(clk), .Q(c2[12]) );
  DFF_X1 c2_reg_11_ ( .D(d[11]), .CK(clk), .Q(c2[11]) );
  DFF_X1 c2_reg_10_ ( .D(d[10]), .CK(clk), .Q(c2[10]) );
  DFF_X1 c2_reg_9_ ( .D(d[9]), .CK(clk), .Q(c2[9]) );
  DFF_X1 c2_reg_8_ ( .D(d[8]), .CK(clk), .Q(c2[8]) );
  DFF_X1 c2_reg_7_ ( .D(d[7]), .CK(clk), .Q(c2[7]) );
  DFF_X1 c2_reg_6_ ( .D(d[6]), .CK(clk), .Q(c2[6]) );
  DFF_X1 c2_reg_5_ ( .D(d[5]), .CK(clk), .Q(c2[5]) );
  DFF_X1 c2_reg_4_ ( .D(d[4]), .CK(clk), .Q(c2[4]) );
  DFF_X1 c2_reg_3_ ( .D(d[3]), .CK(clk), .Q(c2[3]) );
  DFF_X1 c2_reg_2_ ( .D(d[2]), .CK(clk), .Q(c2[2]) );
  DFF_X1 c2_reg_1_ ( .D(d[1]), .CK(clk), .Q(c2[1]) );
  DFF_X1 c2_reg_0_ ( .D(d[0]), .CK(clk), .Q(c2[0]) );
  DFF_X1 c0_reg_17_ ( .D(N464), .CK(clk), .Q(c0[17]) );
  DFF_X1 c0_reg_16_ ( .D(N468), .CK(clk), .Q(c0[16]) );
  DFF_X1 c0_reg_15_ ( .D(N487), .CK(clk), .Q(c0[15]) );
  DFF_X1 c0_reg_14_ ( .D(N509), .CK(clk), .Q(c0[14]) );
  DFF_X1 c0_reg_13_ ( .D(d[48]), .CK(clk), .Q(c0[13]) );
  DFF_X1 c0_reg_12_ ( .D(d[47]), .CK(clk), .Q(c0[12]) );
  DFF_X1 c0_reg_11_ ( .D(d[46]), .CK(clk), .Q(c0[11]) );
  DFF_X1 c0_reg_10_ ( .D(d[45]), .CK(clk), .Q(c0[10]) );
  DFF_X1 c0_reg_9_ ( .D(d[44]), .CK(clk), .Q(c0[9]) );
  DFF_X1 c0_reg_8_ ( .D(d[43]), .CK(clk), .Q(c0[8]) );
  DFF_X1 c0_reg_7_ ( .D(d[42]), .CK(clk), .Q(c0[7]) );
  DFF_X1 c0_reg_6_ ( .D(d[41]), .CK(clk), .Q(c0[6]) );
  DFF_X1 c0_reg_5_ ( .D(d[40]), .CK(clk), .Q(c0[5]) );
  DFF_X1 c0_reg_4_ ( .D(d[39]), .CK(clk), .Q(c0[4]) );
  DFF_X1 c0_reg_3_ ( .D(d[38]), .CK(clk), .Q(c0[3]) );
  DFF_X1 c0_reg_2_ ( .D(d[37]), .CK(clk), .Q(c0[2]) );
  DFF_X1 c0_reg_1_ ( .D(d[36]), .CK(clk), .Q(c0[1]) );
  DFF_X1 c0_reg_0_ ( .D(d[35]), .CK(clk), .Q(c0[0]) );
  DFF_X1 c1_reg_16_ ( .D(N1318), .CK(clk), .Q(c1[16]) );
  DFF_X1 c1_reg_15_ ( .D(N1333), .CK(clk), .Q(c1[15]) );
  DFF_X1 c1_reg_14_ ( .D(N1352), .CK(clk), .Q(c1[14]) );
  DFF_X1 c1_reg_13_ ( .D(d[30]), .CK(clk), .Q(c1[13]) );
  DFF_X1 c1_reg_12_ ( .D(d[29]), .CK(clk), .Q(c1[12]) );
  DFF_X1 c1_reg_11_ ( .D(d[28]), .CK(clk), .Q(c1[11]) );
  DFF_X1 c1_reg_10_ ( .D(d[27]), .CK(clk), .Q(c1[10]) );
  DFF_X1 c1_reg_9_ ( .D(d[26]), .CK(clk), .Q(c1[9]) );
  DFF_X1 c1_reg_8_ ( .D(d[25]), .CK(clk), .Q(c1[8]) );
  DFF_X1 c1_reg_7_ ( .D(d[24]), .CK(clk), .Q(c1[7]) );
  DFF_X1 c1_reg_6_ ( .D(d[23]), .CK(clk), .Q(c1[6]) );
  DFF_X1 c1_reg_5_ ( .D(d[22]), .CK(clk), .Q(c1[5]) );
  DFF_X1 c1_reg_4_ ( .D(d[21]), .CK(clk), .Q(c1[4]) );
  DFF_X1 c1_reg_3_ ( .D(d[20]), .CK(clk), .Q(c1[3]) );
  DFF_X1 c1_reg_2_ ( .D(d[19]), .CK(clk), .Q(c1[2]) );
  DFF_X1 c1_reg_1_ ( .D(d[18]), .CK(clk), .Q(c1[1]) );
  DFF_X1 c1_reg_0_ ( .D(d[17]), .CK(clk), .Q(c1[0]) );
  MUX2_X1 U15 ( .A(n1860), .B(n1857), .S(n1548), .Z(n17) );
  XOR2_X1 U16 ( .A(n473), .B(addr[0]), .Z(n9) );
  MUX2_X1 U19 ( .A(n5), .B(n480), .S(n1548), .Z(n18) );
  MUX2_X1 U21 ( .A(n1857), .B(n463), .S(n1548), .Z(n20) );
  MUX2_X1 U23 ( .A(addr[0]), .B(n2), .S(n1548), .Z(n22) );
  MUX2_X1 U24 ( .A(n444), .B(n2), .S(n1548), .Z(n23) );
  MUX2_X1 U25 ( .A(n1860), .B(addr[0]), .S(n1548), .Z(n24) );
  MUX2_X1 U26 ( .A(n1860), .B(n446), .S(n1548), .Z(n25) );
  MUX2_X1 U27 ( .A(n434), .B(n463), .S(n1548), .Z(n26) );
  XOR2_X1 U29 ( .A(n2), .B(n1544), .Z(n28) );
  MUX2_X1 U31 ( .A(n9), .B(addr[0]), .S(n1548), .Z(n30) );
  MUX2_X1 U32 ( .A(n1858), .B(n463), .S(n1548), .Z(n31) );
  MUX2_X1 U33 ( .A(n1859), .B(n480), .S(n1548), .Z(n32) );
  MUX2_X1 U34 ( .A(n463), .B(n1859), .S(n1548), .Z(n33) );
  MUX2_X1 U35 ( .A(n1858), .B(n480), .S(n1548), .Z(n34) );
  XOR2_X1 U36 ( .A(n1558), .B(n450), .Z(n35) );
  MUX2_X1 U38 ( .A(n1861), .B(n446), .S(n1548), .Z(n37) );
  MUX2_X1 U40 ( .A(addr[0]), .B(n1859), .S(n1548), .Z(n39) );
  MUX2_X1 U41 ( .A(n444), .B(n1861), .S(n1548), .Z(n40) );
  MUX2_X1 U42 ( .A(n1), .B(n5), .S(n1549), .Z(n41) );
  MUX2_X1 U43 ( .A(n1861), .B(n480), .S(n1549), .Z(n42) );
  MUX2_X1 U45 ( .A(n1861), .B(n1859), .S(n1549), .Z(n44) );
  MUX2_X1 U48 ( .A(n9), .B(n1860), .S(n1549), .Z(n47) );
  MUX2_X1 U50 ( .A(n6), .B(n2), .S(n1549), .Z(n49) );
  MUX2_X1 U51 ( .A(n2), .B(addr[0]), .S(n1549), .Z(n50) );
  MUX2_X1 U52 ( .A(n1858), .B(n1861), .S(n1549), .Z(n51) );
  MUX2_X1 U54 ( .A(n2), .B(n1), .S(n1550), .Z(n53) );
  MUX2_X1 U57 ( .A(n1858), .B(n435), .S(n1549), .Z(n56) );
  MUX2_X1 U59 ( .A(n1858), .B(n1859), .S(n1549), .Z(n59) );
  XOR2_X1 U60 ( .A(n506), .B(n1544), .Z(n60) );
  XOR2_X1 U61 ( .A(n498), .B(n450), .Z(n61) );
  XOR2_X1 U62 ( .A(n1558), .B(n1858), .Z(n62) );
  XOR2_X1 U63 ( .A(n4870), .B(n1592), .Z(n63) );
  XOR2_X1 U64 ( .A(n4870), .B(n1859), .Z(n64) );
  XOR2_X1 U65 ( .A(n489), .B(n506), .Z(n65) );
  XOR2_X1 U66 ( .A(n1572), .B(n14), .Z(n66) );
  XOR2_X1 U67 ( .A(n489), .B(n1576), .Z(n67) );
  XOR2_X1 U68 ( .A(n1545), .B(n1576), .Z(n68) );
  XOR2_X1 U69 ( .A(n1559), .B(n1), .Z(n69) );
  MUX2_X1 U70 ( .A(n1645), .B(n1594), .S(n506), .Z(n70) );
  MUX2_X1 U71 ( .A(n1604), .B(n70), .S(n491), .Z(n71) );
  MUX2_X1 U72 ( .A(n1651), .B(n1602), .S(n1520), .Z(n72) );
  MUX2_X1 U73 ( .A(n1652), .B(n1607), .S(n515), .Z(n73) );
  MUX2_X1 U74 ( .A(n73), .B(n72), .S(n493), .Z(n74) );
  MUX2_X1 U75 ( .A(n74), .B(n71), .S(n483), .Z(n75) );
  MUX2_X1 U76 ( .A(addr[0]), .B(n1618), .S(n515), .Z(n76) );
  MUX2_X1 U77 ( .A(n1622), .B(n1620), .S(n515), .Z(n77) );
  MUX2_X1 U78 ( .A(n77), .B(n76), .S(n493), .Z(n78) );
  MUX2_X1 U79 ( .A(n24), .B(n445), .S(n515), .Z(n79) );
  MUX2_X1 U80 ( .A(n1620), .B(n1621), .S(n515), .Z(n80) );
  MUX2_X1 U81 ( .A(n80), .B(n79), .S(n493), .Z(n81) );
  MUX2_X1 U82 ( .A(n81), .B(n78), .S(n484), .Z(n82) );
  MUX2_X1 U83 ( .A(n82), .B(n75), .S(n1576), .Z(n83) );
  MUX2_X1 U84 ( .A(n1619), .B(n1652), .S(n515), .Z(n84) );
  MUX2_X1 U85 ( .A(n1618), .B(addr[0]), .S(n515), .Z(n85) );
  MUX2_X1 U86 ( .A(n85), .B(n84), .S(n493), .Z(n86) );
  MUX2_X1 U87 ( .A(n1857), .B(n446), .S(n515), .Z(n87) );
  MUX2_X1 U88 ( .A(n87), .B(n2), .S(n60), .Z(n88) );
  MUX2_X1 U89 ( .A(n22), .B(n23), .S(n515), .Z(n89) );
  MUX2_X1 U90 ( .A(n89), .B(n88), .S(n493), .Z(n90) );
  MUX2_X1 U91 ( .A(n90), .B(n86), .S(n485), .Z(n91) );
  MUX2_X1 U92 ( .A(n1616), .B(n1617), .S(n515), .Z(n92) );
  MUX2_X1 U93 ( .A(n1614), .B(n1613), .S(n516), .Z(n93) );
  MUX2_X1 U94 ( .A(n93), .B(n92), .S(n493), .Z(n94) );
  MUX2_X1 U95 ( .A(n1653), .B(n3), .S(n516), .Z(n95) );
  MUX2_X1 U96 ( .A(n463), .B(n1858), .S(n1549), .Z(n96) );
  MUX2_X1 U97 ( .A(n1609), .B(n96), .S(n516), .Z(n97) );
  MUX2_X1 U98 ( .A(n97), .B(n95), .S(n493), .Z(n98) );
  MUX2_X1 U99 ( .A(n98), .B(n94), .S(n485), .Z(n99) );
  MUX2_X1 U100 ( .A(n99), .B(n91), .S(n1577), .Z(n100) );
  MUX2_X1 U101 ( .A(n100), .B(n83), .S(n1565), .Z(d[44]) );
  MUX2_X1 U102 ( .A(n1629), .B(n1597), .S(n493), .Z(n101) );
  MUX2_X1 U103 ( .A(n1654), .B(n1596), .S(n493), .Z(n102) );
  MUX2_X1 U104 ( .A(n102), .B(n101), .S(n485), .Z(n103) );
  MUX2_X1 U105 ( .A(n33), .B(n32), .S(n493), .Z(n104) );
  MUX2_X1 U107 ( .A(n105), .B(n8), .S(n493), .Z(n106) );
  MUX2_X1 U108 ( .A(n106), .B(n104), .S(n485), .Z(n107) );
  MUX2_X1 U109 ( .A(n107), .B(n103), .S(n516), .Z(n108) );
  MUX2_X1 U110 ( .A(n34), .B(n33), .S(n493), .Z(n109) );
  MUX2_X1 U111 ( .A(n1858), .B(n1595), .S(n493), .Z(n110) );
  MUX2_X1 U112 ( .A(n110), .B(n109), .S(n485), .Z(n111) );
  MUX2_X1 U113 ( .A(n1627), .B(n1858), .S(n493), .Z(n112) );
  MUX2_X1 U114 ( .A(n1628), .B(n27), .S(n493), .Z(n113) );
  MUX2_X1 U115 ( .A(n113), .B(n112), .S(n485), .Z(n114) );
  MUX2_X1 U116 ( .A(n114), .B(n111), .S(n516), .Z(n115) );
  MUX2_X1 U117 ( .A(n115), .B(n108), .S(addr[7]), .Z(n116) );
  MUX2_X1 U118 ( .A(n5), .B(n6), .S(n1549), .Z(n117) );
  MUX2_X1 U119 ( .A(n9), .B(n117), .S(n493), .Z(n118) );
  MUX2_X1 U120 ( .A(n61), .B(n118), .S(n485), .Z(n119) );
  MUX2_X1 U121 ( .A(n33), .B(n8), .S(n492), .Z(n120) );
  MUX2_X1 U122 ( .A(n1625), .B(n1626), .S(n492), .Z(n121) );
  MUX2_X1 U123 ( .A(n121), .B(n120), .S(n485), .Z(n122) );
  MUX2_X1 U124 ( .A(n122), .B(n119), .S(n516), .Z(n123) );
  MUX2_X1 U125 ( .A(addr[0]), .B(n22), .S(n492), .Z(n124) );
  MUX2_X1 U126 ( .A(n1645), .B(n1651), .S(n492), .Z(n125) );
  MUX2_X1 U127 ( .A(n125), .B(n124), .S(n485), .Z(n126) );
  MUX2_X1 U128 ( .A(n463), .B(n9), .S(n1549), .Z(n127) );
  MUX2_X1 U129 ( .A(n1624), .B(n127), .S(n492), .Z(n128) );
  MUX2_X1 U131 ( .A(n128), .B(n129), .S(n485), .Z(n131) );
  MUX2_X1 U132 ( .A(n131), .B(n126), .S(n516), .Z(n132) );
  MUX2_X1 U133 ( .A(n132), .B(n123), .S(addr[7]), .Z(n133) );
  MUX2_X1 U134 ( .A(n133), .B(n116), .S(n1566), .Z(d[45]) );
  MUX2_X1 U135 ( .A(n1655), .B(n430), .S(n485), .Z(n134) );
  MUX2_X1 U136 ( .A(n134), .B(n1598), .S(n492), .Z(n135) );
  MUX2_X1 U137 ( .A(n12), .B(n411), .S(n492), .Z(n136) );
  MUX2_X1 U138 ( .A(n1562), .B(n136), .S(n429), .Z(n137) );
  MUX2_X1 U139 ( .A(n137), .B(n135), .S(n516), .Z(n138) );
  MUX2_X1 U140 ( .A(n5), .B(n1596), .S(n485), .Z(n139) );
  MUX2_X1 U141 ( .A(n139), .B(n63), .S(n492), .Z(n140) );
  MUX2_X1 U142 ( .A(n1633), .B(n1634), .S(n485), .Z(n141) );
  MUX2_X1 U143 ( .A(n141), .B(n64), .S(n492), .Z(n142) );
  MUX2_X1 U144 ( .A(n142), .B(n140), .S(n516), .Z(n143) );
  MUX2_X1 U145 ( .A(n143), .B(n138), .S(addr[7]), .Z(n144) );
  MUX2_X1 U146 ( .A(n463), .B(n1596), .S(n485), .Z(n145) );
  MUX2_X1 U148 ( .A(n146), .B(n145), .S(n492), .Z(n147) );
  MUX2_X1 U149 ( .A(n32), .B(n5), .S(n485), .Z(n148) );
  MUX2_X1 U150 ( .A(n11), .B(n1597), .S(n485), .Z(n149) );
  MUX2_X1 U151 ( .A(n149), .B(n148), .S(n492), .Z(n150) );
  MUX2_X1 U152 ( .A(n150), .B(n147), .S(n516), .Z(n151) );
  MUX2_X1 U153 ( .A(n1648), .B(n1628), .S(n485), .Z(n152) );
  MUX2_X1 U154 ( .A(n2), .B(n463), .S(n1549), .Z(n153) );
  MUX2_X1 U155 ( .A(n153), .B(n62), .S(n485), .Z(n154) );
  MUX2_X1 U156 ( .A(n154), .B(n152), .S(n492), .Z(n155) );
  MUX2_X1 U157 ( .A(n1631), .B(n1632), .S(n484), .Z(n156) );
  MUX2_X1 U158 ( .A(n1), .B(n463), .S(n1549), .Z(n157) );
  MUX2_X1 U159 ( .A(n157), .B(n1630), .S(n484), .Z(n158) );
  MUX2_X1 U160 ( .A(n158), .B(n156), .S(n492), .Z(n159) );
  MUX2_X1 U161 ( .A(n159), .B(n155), .S(n516), .Z(n160) );
  MUX2_X1 U162 ( .A(n160), .B(n151), .S(addr[7]), .Z(n161) );
  MUX2_X1 U163 ( .A(n161), .B(n144), .S(n1564), .Z(d[46]) );
  MUX2_X1 U164 ( .A(n38), .B(n19), .S(n484), .Z(n162) );
  MUX2_X1 U165 ( .A(n1634), .B(n1552), .S(n484), .Z(n163) );
  MUX2_X1 U166 ( .A(n163), .B(n162), .S(n516), .Z(n164) );
  MUX2_X1 U167 ( .A(n1598), .B(n164), .S(n65), .Z(n165) );
  MUX2_X1 U169 ( .A(n1851), .B(n166), .S(n492), .Z(n167) );
  MUX2_X1 U171 ( .A(n168), .B(n45), .S(n492), .Z(n169) );
  MUX2_X1 U172 ( .A(n169), .B(n167), .S(n516), .Z(n170) );
  MUX2_X1 U173 ( .A(n170), .B(n165), .S(addr[7]), .Z(n171) );
  MUX2_X1 U174 ( .A(n1595), .B(n1552), .S(n484), .Z(n172) );
  MUX2_X1 U175 ( .A(n1561), .B(n172), .S(n492), .Z(n173) );
  MUX2_X1 U176 ( .A(n1552), .B(n411), .S(n484), .Z(n174) );
  MUX2_X1 U177 ( .A(n1557), .B(n12), .S(n484), .Z(n175) );
  MUX2_X1 U178 ( .A(n175), .B(n174), .S(n492), .Z(n176) );
  MUX2_X1 U179 ( .A(n176), .B(n173), .S(n516), .Z(n177) );
  MUX2_X1 U180 ( .A(n1591), .B(n1656), .S(n484), .Z(n178) );
  MUX2_X1 U181 ( .A(n1595), .B(n1635), .S(n484), .Z(n179) );
  MUX2_X1 U182 ( .A(n179), .B(n178), .S(n492), .Z(n180) );
  MUX2_X1 U183 ( .A(n13), .B(n1592), .S(n484), .Z(n181) );
  MUX2_X1 U184 ( .A(n31), .B(n33), .S(n484), .Z(n182) );
  MUX2_X1 U185 ( .A(n182), .B(n181), .S(n491), .Z(n183) );
  MUX2_X1 U186 ( .A(n183), .B(n180), .S(n516), .Z(n184) );
  MUX2_X1 U187 ( .A(n184), .B(n177), .S(addr[7]), .Z(n185) );
  MUX2_X1 U188 ( .A(n185), .B(n171), .S(n1565), .Z(d[47]) );
  MUX2_X1 U189 ( .A(n1636), .B(n1592), .S(n491), .Z(n186) );
  MUX2_X1 U190 ( .A(n14), .B(n186), .S(n1564), .Z(n187) );
  MUX2_X1 U193 ( .A(n189), .B(n188), .S(n1564), .Z(n190) );
  MUX2_X1 U194 ( .A(n190), .B(n187), .S(n484), .Z(n191) );
  MUX2_X1 U195 ( .A(n12), .B(n1552), .S(n491), .Z(n192) );
  MUX2_X1 U197 ( .A(n193), .B(n192), .S(n1564), .Z(n194) );
  MUX2_X1 U198 ( .A(n66), .B(n194), .S(n484), .Z(n195) );
  MUX2_X1 U199 ( .A(n195), .B(n191), .S(n516), .Z(n196) );
  MUX2_X1 U200 ( .A(n12), .B(n427), .S(n491), .Z(n197) );
  MUX2_X1 U202 ( .A(n197), .B(n198), .S(n1564), .Z(n199) );
  MUX2_X1 U204 ( .A(n199), .B(n200), .S(n484), .Z(n202) );
  MUX2_X1 U207 ( .A(n205), .B(n203), .S(n1566), .Z(n206) );
  MUX2_X1 U209 ( .A(n206), .B(n207), .S(n484), .Z(n208) );
  MUX2_X1 U210 ( .A(n208), .B(n202), .S(n516), .Z(n209) );
  MUX2_X1 U211 ( .A(n209), .B(n196), .S(addr[7]), .Z(d[48]) );
  MUX2_X1 U212 ( .A(n1605), .B(n1562), .S(n491), .Z(n210) );
  MUX2_X1 U214 ( .A(n211), .B(n210), .S(n484), .Z(n212) );
  MUX2_X1 U215 ( .A(n105), .B(n1594), .S(n491), .Z(n213) );
  MUX2_X1 U216 ( .A(n427), .B(n1591), .S(n491), .Z(n214) );
  MUX2_X1 U217 ( .A(n214), .B(n213), .S(n484), .Z(n215) );
  MUX2_X1 U218 ( .A(n215), .B(n212), .S(n516), .Z(n216) );
  MUX2_X1 U219 ( .A(n6), .B(n1599), .S(n491), .Z(n217) );
  MUX2_X1 U220 ( .A(n7), .B(n1640), .S(n491), .Z(n218) );
  MUX2_X1 U221 ( .A(n218), .B(n217), .S(n484), .Z(n219) );
  MUX2_X1 U222 ( .A(n221), .B(n1611), .S(n483), .Z(n220) );
  MUX2_X1 U224 ( .A(n222), .B(n219), .S(n1499), .Z(n224) );
  MUX2_X1 U225 ( .A(n224), .B(n216), .S(addr[7]), .Z(n225) );
  MUX2_X1 U226 ( .A(n30), .B(n1639), .S(n491), .Z(n226) );
  MUX2_X1 U227 ( .A(n411), .B(n1638), .S(n491), .Z(n227) );
  MUX2_X1 U228 ( .A(n227), .B(n226), .S(n483), .Z(n228) );
  MUX2_X1 U229 ( .A(n26), .B(n39), .S(n491), .Z(n229) );
  MUX2_X1 U230 ( .A(n37), .B(n15), .S(n491), .Z(n230) );
  MUX2_X1 U231 ( .A(n230), .B(n229), .S(n483), .Z(n231) );
  MUX2_X1 U232 ( .A(n231), .B(n228), .S(n1499), .Z(n232) );
  MUX2_X1 U233 ( .A(n1611), .B(n445), .S(n491), .Z(n233) );
  MUX2_X1 U234 ( .A(n233), .B(n1597), .S(n483), .Z(n234) );
  MUX2_X1 U235 ( .A(n1857), .B(n1859), .S(n1549), .Z(n235) );
  MUX2_X1 U236 ( .A(n2), .B(n6), .S(n1549), .Z(n236) );
  MUX2_X1 U237 ( .A(n236), .B(n235), .S(n491), .Z(n237) );
  MUX2_X1 U238 ( .A(n1631), .B(n1637), .S(n491), .Z(n238) );
  MUX2_X1 U239 ( .A(n238), .B(n237), .S(n483), .Z(n239) );
  MUX2_X1 U240 ( .A(n239), .B(n234), .S(n1499), .Z(n240) );
  MUX2_X1 U241 ( .A(n240), .B(n232), .S(addr[7]), .Z(n241) );
  MUX2_X1 U242 ( .A(n241), .B(n225), .S(n1564), .Z(d[4]) );
  MUX2_X1 U243 ( .A(n1606), .B(n1591), .S(n1578), .Z(n242) );
  MUX2_X1 U244 ( .A(n478), .B(n1859), .S(n1549), .Z(n243) );
  MUX2_X1 U245 ( .A(n243), .B(n1605), .S(addr[7]), .Z(n244) );
  MUX2_X1 U246 ( .A(n244), .B(n242), .S(n491), .Z(n245) );
  MUX2_X1 U247 ( .A(n1650), .B(n1597), .S(n1579), .Z(n246) );
  MUX2_X1 U249 ( .A(n247), .B(n246), .S(n491), .Z(n249) );
  MUX2_X1 U250 ( .A(n249), .B(n245), .S(n483), .Z(n250) );
  MUX2_X1 U251 ( .A(n1615), .B(n1592), .S(n1577), .Z(n251) );
  MUX2_X1 U253 ( .A(n252), .B(n251), .S(n490), .Z(n253) );
  MUX2_X1 U254 ( .A(n43), .B(n1640), .S(n490), .Z(n254) );
  MUX2_X1 U255 ( .A(n254), .B(n1655), .S(n67), .Z(n255) );
  MUX2_X1 U256 ( .A(n255), .B(n253), .S(n483), .Z(n256) );
  MUX2_X1 U257 ( .A(n256), .B(n250), .S(n1499), .Z(n257) );
  MUX2_X1 U258 ( .A(n1656), .B(n1657), .S(addr[7]), .Z(n258) );
  MUX2_X1 U260 ( .A(n258), .B(n259), .S(n490), .Z(n260) );
  MUX2_X1 U263 ( .A(n58), .B(n261), .S(addr[7]), .Z(n262) );
  MUX2_X1 U264 ( .A(n47), .B(n1), .S(addr[7]), .Z(n263) );
  MUX2_X1 U265 ( .A(n263), .B(n262), .S(n490), .Z(n264) );
  MUX2_X1 U266 ( .A(n264), .B(n260), .S(n483), .Z(n265) );
  MUX2_X1 U267 ( .A(n1658), .B(n26), .S(addr[7]), .Z(n266) );
  MUX2_X1 U269 ( .A(n267), .B(n266), .S(n490), .Z(n268) );
  MUX2_X1 U270 ( .A(n5), .B(n1860), .S(n1579), .Z(n269) );
  MUX2_X1 U271 ( .A(n269), .B(n1859), .S(n68), .Z(n270) );
  MUX2_X1 U272 ( .A(n477), .B(n1860), .S(n1549), .Z(n271) );
  MUX2_X1 U273 ( .A(n27), .B(n271), .S(n1579), .Z(n272) );
  MUX2_X1 U274 ( .A(n272), .B(n270), .S(n490), .Z(n273) );
  MUX2_X1 U275 ( .A(n273), .B(n268), .S(n483), .Z(n274) );
  MUX2_X1 U276 ( .A(n274), .B(n265), .S(n1499), .Z(n275) );
  MUX2_X1 U277 ( .A(n275), .B(n257), .S(n1564), .Z(d[5]) );
  MUX2_X1 U278 ( .A(n1591), .B(n1592), .S(n483), .Z(n276) );
  MUX2_X1 U279 ( .A(n1600), .B(n276), .S(n429), .Z(n277) );
  MUX2_X1 U280 ( .A(n1647), .B(n1594), .S(n490), .Z(n278) );
  MUX2_X1 U281 ( .A(n1625), .B(n1629), .S(n490), .Z(n279) );
  MUX2_X1 U282 ( .A(n279), .B(n278), .S(n483), .Z(n280) );
  MUX2_X1 U283 ( .A(n280), .B(n277), .S(n1499), .Z(n281) );
  MUX2_X1 U284 ( .A(n1594), .B(n1622), .S(n490), .Z(n282) );
  MUX2_X1 U285 ( .A(n1659), .B(n40), .S(n490), .Z(n283) );
  MUX2_X1 U286 ( .A(n283), .B(n282), .S(n483), .Z(n284) );
  MUX2_X1 U287 ( .A(n21), .B(n4), .S(n490), .Z(n285) );
  MUX2_X1 U288 ( .A(n1633), .B(n1641), .S(n490), .Z(n286) );
  MUX2_X1 U289 ( .A(n286), .B(n285), .S(n483), .Z(n287) );
  MUX2_X1 U290 ( .A(n287), .B(n284), .S(n1499), .Z(n288) );
  MUX2_X1 U291 ( .A(n288), .B(n281), .S(n1579), .Z(n289) );
  MUX2_X1 U292 ( .A(n1660), .B(n53), .S(n490), .Z(n290) );
  MUX2_X1 U293 ( .A(n15), .B(n1640), .S(n490), .Z(n291) );
  MUX2_X1 U294 ( .A(n291), .B(n290), .S(n483), .Z(n292) );
  MUX2_X1 U295 ( .A(n1637), .B(n16), .S(n490), .Z(n293) );
  MUX2_X1 U296 ( .A(n50), .B(n35), .S(n490), .Z(n294) );
  MUX2_X1 U297 ( .A(n294), .B(n293), .S(n483), .Z(n295) );
  MUX2_X1 U298 ( .A(n295), .B(n292), .S(n1499), .Z(n296) );
  MUX2_X1 U299 ( .A(n1610), .B(n54), .S(n490), .Z(n297) );
  MUX2_X1 U301 ( .A(n298), .B(n297), .S(n483), .Z(n299) );
  MUX2_X1 U302 ( .A(n1660), .B(n1641), .S(n490), .Z(n300) );
  MUX2_X1 U303 ( .A(n1612), .B(n1661), .S(n492), .Z(n301) );
  MUX2_X1 U304 ( .A(n301), .B(n300), .S(n483), .Z(n302) );
  MUX2_X1 U305 ( .A(n302), .B(n299), .S(n1499), .Z(n303) );
  MUX2_X1 U306 ( .A(n303), .B(n296), .S(n1579), .Z(n304) );
  MUX2_X1 U307 ( .A(n304), .B(n289), .S(n1565), .Z(d[6]) );
  MUX2_X1 U308 ( .A(n1599), .B(n1562), .S(n490), .Z(n305) );
  MUX2_X1 U310 ( .A(n306), .B(n305), .S(n482), .Z(n307) );
  MUX2_X1 U311 ( .A(n1860), .B(n9), .S(n1550), .Z(n308) );
  MUX2_X1 U312 ( .A(n1626), .B(n308), .S(n490), .Z(n309) );
  MUX2_X1 U314 ( .A(n309), .B(n310), .S(n482), .Z(n312) );
  MUX2_X1 U315 ( .A(n312), .B(n307), .S(n1499), .Z(n313) );
  MUX2_X1 U316 ( .A(n444), .B(n1), .S(n1550), .Z(n314) );
  MUX2_X1 U317 ( .A(n314), .B(n1595), .S(n492), .Z(n315) );
  MUX2_X1 U319 ( .A(n315), .B(n316), .S(n482), .Z(n318) );
  MUX2_X1 U320 ( .A(n25), .B(n51), .S(n491), .Z(n319) );
  MUX2_X1 U321 ( .A(n5), .B(addr[0]), .S(n1550), .Z(n320) );
  MUX2_X1 U322 ( .A(n444), .B(n320), .S(n489), .Z(n321) );
  MUX2_X1 U323 ( .A(n321), .B(n319), .S(n482), .Z(n322) );
  MUX2_X1 U324 ( .A(n322), .B(n318), .S(n1499), .Z(n323) );
  MUX2_X1 U325 ( .A(n323), .B(n313), .S(n1579), .Z(n324) );
  MUX2_X1 U326 ( .A(n1653), .B(n1562), .S(n491), .Z(n325) );
  MUX2_X1 U327 ( .A(n1639), .B(n8), .S(n492), .Z(n326) );
  MUX2_X1 U328 ( .A(n326), .B(n325), .S(n482), .Z(n327) );
  MUX2_X1 U330 ( .A(n328), .B(n7), .S(n490), .Z(n329) );
  MUX2_X1 U331 ( .A(n1625), .B(n1612), .S(n491), .Z(n330) );
  MUX2_X1 U332 ( .A(n330), .B(n329), .S(n482), .Z(n331) );
  MUX2_X1 U333 ( .A(n331), .B(n327), .S(n1499), .Z(n332) );
  MUX2_X1 U334 ( .A(n1634), .B(n1625), .S(n491), .Z(n333) );
  MUX2_X1 U335 ( .A(n56), .B(n1608), .S(n489), .Z(n334) );
  MUX2_X1 U336 ( .A(n334), .B(n333), .S(n482), .Z(n335) );
  MUX2_X1 U337 ( .A(n1599), .B(n5), .S(n489), .Z(n336) );
  MUX2_X1 U338 ( .A(n1603), .B(n31), .S(n489), .Z(n337) );
  MUX2_X1 U339 ( .A(n337), .B(n336), .S(n482), .Z(n338) );
  MUX2_X1 U340 ( .A(n338), .B(n335), .S(n1499), .Z(n339) );
  MUX2_X1 U341 ( .A(n339), .B(n332), .S(n1579), .Z(n340) );
  MUX2_X1 U342 ( .A(n340), .B(n324), .S(n1566), .Z(d[7]) );
  MUX2_X1 U343 ( .A(n430), .B(n69), .S(n489), .Z(n341) );
  MUX2_X1 U345 ( .A(n56), .B(n342), .S(n1579), .Z(n343) );
  MUX2_X1 U346 ( .A(n1605), .B(n1599), .S(n1579), .Z(n344) );
  MUX2_X1 U347 ( .A(n344), .B(n343), .S(n489), .Z(n345) );
  MUX2_X1 U349 ( .A(n345), .B(n346), .S(n482), .Z(n348) );
  MUX2_X1 U350 ( .A(n5), .B(n9), .S(n1550), .Z(n349) );
  MUX2_X1 U351 ( .A(n52), .B(n349), .S(n1579), .Z(n350) );
  MUX2_X1 U353 ( .A(n350), .B(n351), .S(n489), .Z(n352) );
  MUX2_X1 U354 ( .A(n1638), .B(n1607), .S(n1579), .Z(n353) );
  MUX2_X1 U356 ( .A(n353), .B(n354), .S(n489), .Z(n355) );
  MUX2_X1 U357 ( .A(n355), .B(n352), .S(n482), .Z(n356) );
  MUX2_X1 U358 ( .A(n356), .B(n348), .S(n1499), .Z(n357) );
  MUX2_X1 U360 ( .A(n36), .B(n358), .S(n1579), .Z(n359) );
  MUX2_X1 U361 ( .A(n41), .B(n20), .S(n1579), .Z(n360) );
  MUX2_X1 U362 ( .A(n360), .B(n359), .S(n489), .Z(n361) );
  MUX2_X1 U363 ( .A(n3), .B(n1622), .S(n1579), .Z(n362) );
  MUX2_X1 U364 ( .A(n6), .B(n1), .S(n1550), .Z(n363) );
  MUX2_X1 U365 ( .A(n363), .B(n12), .S(n1579), .Z(n364) );
  MUX2_X1 U366 ( .A(n364), .B(n362), .S(n493), .Z(n365) );
  MUX2_X1 U367 ( .A(n365), .B(n361), .S(n482), .Z(n366) );
  MUX2_X1 U368 ( .A(n1617), .B(n19), .S(n1579), .Z(n367) );
  MUX2_X1 U369 ( .A(n9), .B(n46), .S(n1579), .Z(n368) );
  MUX2_X1 U370 ( .A(n368), .B(n367), .S(n489), .Z(n369) );
  MUX2_X1 U371 ( .A(n463), .B(n1658), .S(n1579), .Z(n370) );
  MUX2_X1 U372 ( .A(addr[0]), .B(n1861), .S(n1550), .Z(n371) );
  MUX2_X1 U373 ( .A(n16), .B(n371), .S(n1579), .Z(n372) );
  MUX2_X1 U374 ( .A(n372), .B(n370), .S(n489), .Z(n373) );
  MUX2_X1 U375 ( .A(n373), .B(n369), .S(n482), .Z(n374) );
  MUX2_X1 U376 ( .A(n374), .B(n366), .S(n1499), .Z(n375) );
  MUX2_X1 U377 ( .A(n375), .B(n357), .S(n1566), .Z(d[8]) );
  MUX2_X1 U378 ( .A(n1597), .B(n1593), .S(n1499), .Z(n376) );
  MUX2_X1 U379 ( .A(n1604), .B(n376), .S(n489), .Z(n377) );
  MUX2_X1 U380 ( .A(n1595), .B(n1592), .S(n1499), .Z(n378) );
  MUX2_X1 U382 ( .A(n379), .B(n378), .S(n489), .Z(n380) );
  MUX2_X1 U383 ( .A(n380), .B(n377), .S(n482), .Z(n381) );
  MUX2_X1 U384 ( .A(n49), .B(n1631), .S(n1499), .Z(n382) );
  MUX2_X1 U385 ( .A(n1616), .B(n1659), .S(n1500), .Z(n383) );
  MUX2_X1 U386 ( .A(n383), .B(n382), .S(n489), .Z(n384) );
  MUX2_X1 U387 ( .A(n1592), .B(n1649), .S(n1500), .Z(n385) );
  MUX2_X1 U388 ( .A(n57), .B(n1642), .S(n1500), .Z(n386) );
  MUX2_X1 U389 ( .A(n386), .B(n385), .S(n492), .Z(n387) );
  MUX2_X1 U390 ( .A(n387), .B(n384), .S(n482), .Z(n388) );
  MUX2_X1 U391 ( .A(n388), .B(n381), .S(n1579), .Z(n389) );
  MUX2_X1 U392 ( .A(n1662), .B(n1638), .S(n1500), .Z(n390) );
  MUX2_X1 U393 ( .A(n55), .B(n59), .S(n1500), .Z(n391) );
  MUX2_X1 U394 ( .A(n391), .B(n390), .S(n489), .Z(n392) );
  MUX2_X1 U395 ( .A(n52), .B(n1657), .S(n1500), .Z(n393) );
  MUX2_X1 U396 ( .A(n444), .B(n1859), .S(n1550), .Z(n394) );
  MUX2_X1 U397 ( .A(n1654), .B(n394), .S(n1500), .Z(n395) );
  MUX2_X1 U398 ( .A(n395), .B(n393), .S(n490), .Z(n396) );
  MUX2_X1 U399 ( .A(n396), .B(n392), .S(n482), .Z(n397) );
  MUX2_X1 U400 ( .A(n41), .B(n1662), .S(n1500), .Z(n398) );
  MUX2_X1 U401 ( .A(n1), .B(n1644), .S(n1500), .Z(n399) );
  MUX2_X1 U402 ( .A(n399), .B(n398), .S(n489), .Z(n400) );
  MUX2_X1 U404 ( .A(n400), .B(n401), .S(n482), .Z(n404) );
  MUX2_X1 U405 ( .A(n404), .B(n397), .S(n1578), .Z(n405) );
  MUX2_X1 U406 ( .A(n405), .B(n389), .S(n1564), .Z(d[9]) );
  MUX2_X1 U407 ( .A(n9), .B(n1857), .S(n1550), .Z(n221) );
  MUX2_X1 U420 ( .A(n1623), .B(n407), .S(n1500), .Z(n412) );
  MUX2_X1 U421 ( .A(n444), .B(n9), .S(n1550), .Z(n413) );
  MUX2_X1 U422 ( .A(n2), .B(n1858), .S(n1550), .Z(n414) );
  MUX2_X1 U423 ( .A(n1860), .B(n463), .S(n1550), .Z(n415) );
  MUX2_X1 U424 ( .A(n476), .B(n6), .S(n1550), .Z(n416) );
  MUX2_X1 U425 ( .A(n1552), .B(n38), .S(n482), .Z(n417) );
  MUX2_X1 U426 ( .A(n475), .B(n1861), .S(n1550), .Z(n418) );
  MUX2_X1 U427 ( .A(n1861), .B(n463), .S(n1550), .Z(n419) );
  MUX2_X1 U428 ( .A(n1646), .B(n1562), .S(n489), .Z(n201) );
  MUX2_X1 U429 ( .A(n41), .B(n43), .S(n482), .Z(n223) );
  MUX2_X1 U430 ( .A(n463), .B(n2), .S(n1550), .Z(n420) );
  MUX2_X1 U431 ( .A(n5), .B(n2), .S(n1550), .Z(n421) );
  MUX2_X1 U432 ( .A(n1861), .B(n1858), .S(n1551), .Z(n422) );
  MUX2_X1 U433 ( .A(n473), .B(n1), .S(n1550), .Z(n423) );
  MUX2_X1 U434 ( .A(addr[0]), .B(n1), .S(n1551), .Z(n424) );
  MUX2_X1 U435 ( .A(n406), .B(n13), .S(n490), .Z(n347) );
  MUX2_X1 U436 ( .A(addr[0]), .B(n9), .S(n1551), .Z(n425) );
  MUX2_X1 U438 ( .A(n426), .B(n1525), .S(n489), .Z(n403) );
  MUX2_X1 U439 ( .A(n1614), .B(n1610), .S(n489), .Z(n402) );
  XOR2_X1 U554 ( .A(n498), .B(addr[2]), .Z(n533) );
  MUX2_X1 U556 ( .A(n4870), .B(n1829), .S(n435), .Z(n549) );
  MUX2_X1 U557 ( .A(n1843), .B(n533), .S(n435), .Z(n550) );
  MUX2_X1 U563 ( .A(n1829), .B(n1750), .S(n435), .Z(n553) );
  MUX2_X1 U564 ( .A(n501), .B(n1782), .S(n435), .Z(n554) );
  MUX2_X1 U566 ( .A(n528), .B(n520), .S(n435), .Z(n556) );
  MUX2_X1 U567 ( .A(n533), .B(n492), .S(n435), .Z(n557) );
  MUX2_X1 U569 ( .A(n528), .B(n517), .S(n435), .Z(n559) );
  XOR2_X1 U571 ( .A(n440), .B(n1782), .Z(n561) );
  MUX2_X1 U572 ( .A(n493), .B(n483), .S(n434), .Z(n562) );
  MUX2_X1 U573 ( .A(n1782), .B(n517), .S(n435), .Z(n563) );
  MUX2_X1 U574 ( .A(n483), .B(n1782), .S(n435), .Z(n564) );
  MUX2_X1 U575 ( .A(n533), .B(n526), .S(n435), .Z(n565) );
  MUX2_X1 U576 ( .A(n1800), .B(n1829), .S(n435), .Z(n566) );
  MUX2_X1 U577 ( .A(n501), .B(n526), .S(n435), .Z(n567) );
  XOR2_X1 U578 ( .A(n1559), .B(n506), .Z(n568) );
  MUX2_X1 U580 ( .A(n483), .B(n528), .S(n435), .Z(n570) );
  MUX2_X1 U581 ( .A(n1782), .B(n492), .S(n435), .Z(n571) );
  MUX2_X1 U582 ( .A(n1843), .B(n1800), .S(n435), .Z(n572) );
  MUX2_X1 U583 ( .A(n493), .B(n520), .S(n435), .Z(n547) );
  MUX2_X1 U584 ( .A(n501), .B(n533), .S(n434), .Z(n573) );
  MUX2_X1 U586 ( .A(n517), .B(n483), .S(n434), .Z(n575) );
  MUX2_X1 U587 ( .A(n482), .B(n1843), .S(n434), .Z(n576) );
  MUX2_X1 U588 ( .A(n520), .B(n526), .S(n434), .Z(n577) );
  MUX2_X1 U589 ( .A(n520), .B(n492), .S(n434), .Z(n578) );
  XOR2_X1 U590 ( .A(n499), .B(n432), .Z(n579) );
  MUX2_X1 U594 ( .A(n533), .B(n483), .S(n434), .Z(n583) );
  MUX2_X1 U595 ( .A(n1750), .B(n484), .S(n434), .Z(n584) );
  MUX2_X1 U596 ( .A(n1750), .B(n1800), .S(n434), .Z(n585) );
  MUX2_X1 U597 ( .A(n517), .B(n502), .S(n434), .Z(n586) );
  MUX2_X1 U599 ( .A(n493), .B(n526), .S(n434), .Z(n588) );
  MUX2_X1 U600 ( .A(n483), .B(n1800), .S(n434), .Z(n589) );
  XOR2_X1 U601 ( .A(n517), .B(n432), .Z(n590) );
  MUX2_X1 U602 ( .A(n1829), .B(n1782), .S(n434), .Z(n591) );
  MUX2_X1 U605 ( .A(n4870), .B(n517), .S(n434), .Z(n594) );
  MUX2_X1 U606 ( .A(n526), .B(n484), .S(n434), .Z(n595) );
  MUX2_X1 U607 ( .A(n1829), .B(n482), .S(n434), .Z(n596) );
  MUX2_X1 U609 ( .A(n485), .B(n489), .S(n434), .Z(n598) );
  MUX2_X1 U610 ( .A(n500), .B(n528), .S(n434), .Z(n599) );
  MUX2_X1 U612 ( .A(n1800), .B(n501), .S(n433), .Z(n601) );
  MUX2_X1 U613 ( .A(n499), .B(n483), .S(n433), .Z(n602) );
  MUX2_X1 U614 ( .A(n517), .B(n1782), .S(n433), .Z(n603) );
  MUX2_X1 U616 ( .A(n1800), .B(n1782), .S(n433), .Z(n605) );
  MUX2_X1 U617 ( .A(n1782), .B(n484), .S(n433), .Z(n606) );
  MUX2_X1 U619 ( .A(n533), .B(n1843), .S(n433), .Z(n608) );
  MUX2_X1 U620 ( .A(n1750), .B(n1843), .S(n433), .Z(n609) );
  MUX2_X1 U621 ( .A(n533), .B(n520), .S(n433), .Z(n610) );
  MUX2_X1 U622 ( .A(n520), .B(n528), .S(n433), .Z(n611) );
  MUX2_X1 U623 ( .A(n526), .B(n502), .S(n433), .Z(n612) );
  MUX2_X1 U624 ( .A(n528), .B(n482), .S(n433), .Z(n613) );
  MUX2_X1 U625 ( .A(n1829), .B(n4870), .S(n433), .Z(n614) );
  MUX2_X1 U626 ( .A(n4870), .B(n1782), .S(n433), .Z(n615) );
  MUX2_X1 U628 ( .A(n4870), .B(n1750), .S(n433), .Z(n617) );
  MUX2_X1 U629 ( .A(n496), .B(n1750), .S(n433), .Z(n618) );
  MUX2_X1 U630 ( .A(n489), .B(n1829), .S(n433), .Z(n619) );
  MUX2_X1 U631 ( .A(n1843), .B(n484), .S(n432), .Z(n620) );
  MUX2_X1 U632 ( .A(n1750), .B(n501), .S(n433), .Z(n621) );
  MUX2_X1 U633 ( .A(n1829), .B(n490), .S(n432), .Z(n622) );
  MUX2_X1 U634 ( .A(n443), .B(n1792), .S(n1500), .Z(n623) );
  XOR2_X1 U637 ( .A(n528), .B(n432), .Z(n626) );
  XOR2_X1 U638 ( .A(n526), .B(n433), .Z(n627) );
  XOR2_X1 U639 ( .A(n520), .B(n432), .Z(n628) );
  XOR2_X1 U640 ( .A(n4870), .B(n433), .Z(n629) );
  XOR2_X1 U641 ( .A(n539), .B(n506), .Z(n630) );
  XOR2_X1 U642 ( .A(n1534), .B(n1809), .Z(n631) );
  XOR2_X1 U643 ( .A(n1534), .B(n432), .Z(n632) );
  XOR2_X1 U644 ( .A(n517), .B(n506), .Z(n633) );
  MUX2_X1 U645 ( .A(n1808), .B(n1765), .S(n1568), .Z(n634) );
  MUX2_X1 U647 ( .A(n634), .B(n635), .S(n1500), .Z(n636) );
  MUX2_X1 U648 ( .A(n1773), .B(n1789), .S(addr[6]), .Z(n637) );
  MUX2_X1 U650 ( .A(n637), .B(n638), .S(n1500), .Z(n639) );
  MUX2_X1 U651 ( .A(n639), .B(n636), .S(n457), .Z(n640) );
  MUX2_X1 U652 ( .A(n550), .B(n530), .S(n1568), .Z(n641) );
  MUX2_X1 U653 ( .A(n521), .B(n1835), .S(n1568), .Z(n642) );
  MUX2_X1 U654 ( .A(n642), .B(n641), .S(n1500), .Z(n643) );
  MUX2_X1 U655 ( .A(n1855), .B(addr[0]), .S(addr[6]), .Z(n644) );
  MUX2_X1 U656 ( .A(n1674), .B(n1772), .S(addr[6]), .Z(n645) );
  MUX2_X1 U657 ( .A(n645), .B(n644), .S(n1500), .Z(n646) );
  MUX2_X1 U658 ( .A(n646), .B(n643), .S(n457), .Z(n647) );
  MUX2_X1 U659 ( .A(n647), .B(n640), .S(n1551), .Z(n648) );
  MUX2_X1 U660 ( .A(n1792), .B(n1754), .S(n1568), .Z(n649) );
  MUX2_X1 U661 ( .A(n526), .B(n1823), .S(addr[6]), .Z(n650) );
  MUX2_X1 U662 ( .A(n650), .B(n649), .S(n1500), .Z(n651) );
  MUX2_X1 U663 ( .A(n527), .B(n529), .S(addr[6]), .Z(n652) );
  MUX2_X1 U664 ( .A(n628), .B(n524), .S(addr[6]), .Z(n653) );
  MUX2_X1 U665 ( .A(n653), .B(n652), .S(n1500), .Z(n654) );
  MUX2_X1 U666 ( .A(n654), .B(n651), .S(n457), .Z(n655) );
  MUX2_X1 U667 ( .A(n1800), .B(n1792), .S(addr[6]), .Z(n656) );
  MUX2_X1 U668 ( .A(n1822), .B(n1790), .S(addr[6]), .Z(n657) );
  MUX2_X1 U669 ( .A(n657), .B(n656), .S(n1500), .Z(n658) );
  MUX2_X1 U670 ( .A(n518), .B(n1769), .S(n1568), .Z(n659) );
  MUX2_X1 U672 ( .A(n659), .B(n660), .S(n1501), .Z(n661) );
  MUX2_X1 U673 ( .A(n661), .B(n658), .S(n457), .Z(n662) );
  MUX2_X1 U674 ( .A(n662), .B(n655), .S(n1551), .Z(n663) );
  MUX2_X1 U675 ( .A(n663), .B(n648), .S(n1578), .Z(d[0]) );
  MUX2_X1 U676 ( .A(n1793), .B(n1829), .S(n1551), .Z(n664) );
  MUX2_X1 U678 ( .A(n665), .B(n1663), .S(n457), .Z(n666) );
  MUX2_X1 U679 ( .A(n536), .B(addr[0]), .S(n1501), .Z(n667) );
  MUX2_X1 U680 ( .A(n534), .B(n667), .S(n1551), .Z(n668) );
  MUX2_X1 U681 ( .A(n1802), .B(n524), .S(n1501), .Z(n669) );
  MUX2_X1 U682 ( .A(n532), .B(n1807), .S(n1501), .Z(n670) );
  MUX2_X1 U683 ( .A(n670), .B(n669), .S(n1551), .Z(n671) );
  MUX2_X1 U684 ( .A(n671), .B(n668), .S(n457), .Z(n672) );
  MUX2_X1 U685 ( .A(n672), .B(n666), .S(n1565), .Z(n673) );
  MUX2_X1 U686 ( .A(n1829), .B(n535), .S(n1501), .Z(n674) );
  MUX2_X1 U688 ( .A(n675), .B(n674), .S(n1551), .Z(n676) );
  MUX2_X1 U689 ( .A(n1788), .B(n1789), .S(n1501), .Z(n677) );
  MUX2_X1 U690 ( .A(n629), .B(n533), .S(n1501), .Z(n678) );
  MUX2_X1 U691 ( .A(n678), .B(n677), .S(n1551), .Z(n679) );
  MUX2_X1 U692 ( .A(n679), .B(n676), .S(n457), .Z(n680) );
  MUX2_X1 U693 ( .A(n1764), .B(n1775), .S(n1501), .Z(n681) );
  MUX2_X1 U694 ( .A(n1811), .B(n1820), .S(n1501), .Z(n682) );
  MUX2_X1 U695 ( .A(n682), .B(n681), .S(n1551), .Z(n683) );
  MUX2_X1 U696 ( .A(n522), .B(n1848), .S(n1501), .Z(n684) );
  MUX2_X1 U697 ( .A(n517), .B(n1774), .S(n1501), .Z(n685) );
  MUX2_X1 U698 ( .A(n685), .B(n684), .S(n1551), .Z(n686) );
  MUX2_X1 U699 ( .A(n686), .B(n683), .S(n458), .Z(n687) );
  MUX2_X1 U700 ( .A(n687), .B(n680), .S(n1568), .Z(n688) );
  MUX2_X1 U701 ( .A(n688), .B(n673), .S(n1578), .Z(d[10]) );
  MUX2_X1 U703 ( .A(n689), .B(n1665), .S(n1551), .Z(n690) );
  MUX2_X1 U704 ( .A(n690), .B(n1663), .S(n458), .Z(n691) );
  MUX2_X1 U706 ( .A(n1670), .B(n692), .S(n1551), .Z(n693) );
  MUX2_X1 U708 ( .A(n693), .B(n694), .S(n458), .Z(n695) );
  MUX2_X1 U709 ( .A(n695), .B(n691), .S(n1568), .Z(n696) );
  MUX2_X1 U710 ( .A(n630), .B(n574), .S(n1551), .Z(n697) );
  MUX2_X1 U711 ( .A(n1787), .B(n1829), .S(n1501), .Z(n698) );
  MUX2_X1 U712 ( .A(n698), .B(n631), .S(n1551), .Z(n699) );
  MUX2_X1 U713 ( .A(n699), .B(n697), .S(n458), .Z(n700) );
  MUX2_X1 U714 ( .A(n1796), .B(n1833), .S(n1501), .Z(n701) );
  MUX2_X1 U715 ( .A(n1837), .B(n4870), .S(n1501), .Z(n702) );
  MUX2_X1 U716 ( .A(n702), .B(n701), .S(n1551), .Z(n703) );
  MUX2_X1 U717 ( .A(n1846), .B(n1776), .S(n1501), .Z(n704) );
  MUX2_X1 U718 ( .A(n604), .B(n538), .S(n1501), .Z(n705) );
  MUX2_X1 U719 ( .A(n705), .B(n704), .S(n1552), .Z(n706) );
  MUX2_X1 U720 ( .A(n706), .B(n703), .S(n458), .Z(n707) );
  MUX2_X1 U721 ( .A(n707), .B(n700), .S(n1568), .Z(n708) );
  MUX2_X1 U722 ( .A(n708), .B(n696), .S(n1578), .Z(d[11]) );
  MUX2_X1 U723 ( .A(n1792), .B(n537), .S(n1568), .Z(n709) );
  MUX2_X1 U725 ( .A(n710), .B(n709), .S(n1501), .Z(n711) );
  MUX2_X1 U727 ( .A(n711), .B(n712), .S(n1549), .Z(n713) );
  MUX2_X1 U729 ( .A(n713), .B(n714), .S(n458), .Z(n715) );
  MUX2_X1 U730 ( .A(n531), .B(n445), .S(n1568), .Z(n716) );
  MUX2_X1 U732 ( .A(n717), .B(n716), .S(n1501), .Z(n718) );
  MUX2_X1 U733 ( .A(n489), .B(addr[0]), .S(n1568), .Z(n719) );
  MUX2_X1 U734 ( .A(n569), .B(n536), .S(n1568), .Z(n720) );
  MUX2_X1 U735 ( .A(n720), .B(n719), .S(n1520), .Z(n721) );
  MUX2_X1 U736 ( .A(n721), .B(n718), .S(n1544), .Z(n722) );
  MUX2_X1 U737 ( .A(n535), .B(n539), .S(n1568), .Z(n723) );
  MUX2_X1 U738 ( .A(n495), .B(addr[0]), .S(n1568), .Z(n724) );
  MUX2_X1 U739 ( .A(n724), .B(n723), .S(n1520), .Z(n725) );
  MUX2_X1 U740 ( .A(n1839), .B(n628), .S(n1568), .Z(n726) );
  MUX2_X1 U741 ( .A(n1763), .B(n1807), .S(n1568), .Z(n727) );
  MUX2_X1 U742 ( .A(n727), .B(n726), .S(n1520), .Z(n728) );
  MUX2_X1 U743 ( .A(n728), .B(n725), .S(n1546), .Z(n729) );
  MUX2_X1 U744 ( .A(n729), .B(n722), .S(n458), .Z(n730) );
  MUX2_X1 U745 ( .A(n730), .B(n715), .S(n1578), .Z(d[12]) );
  MUX2_X1 U746 ( .A(n531), .B(n1829), .S(n458), .Z(n731) );
  MUX2_X1 U749 ( .A(n733), .B(n732), .S(n1545), .Z(n735) );
  MUX2_X1 U751 ( .A(n736), .B(n735), .S(n1568), .Z(n737) );
  MUX2_X1 U752 ( .A(n581), .B(n1837), .S(n1520), .Z(n738) );
  MUX2_X1 U753 ( .A(n738), .B(addr[0]), .S(n458), .Z(n739) );
  MUX2_X1 U755 ( .A(n739), .B(n740), .S(n1547), .Z(n741) );
  MUX2_X1 U758 ( .A(n743), .B(n742), .S(n1520), .Z(n744) );
  MUX2_X1 U759 ( .A(n547), .B(n1812), .S(n458), .Z(n745) );
  MUX2_X1 U760 ( .A(n1832), .B(n577), .S(n458), .Z(n746) );
  MUX2_X1 U761 ( .A(n746), .B(n745), .S(n1520), .Z(n747) );
  MUX2_X1 U762 ( .A(n747), .B(n744), .S(n1546), .Z(n748) );
  MUX2_X1 U763 ( .A(n748), .B(n741), .S(n1568), .Z(n749) );
  MUX2_X1 U764 ( .A(n749), .B(n737), .S(n1578), .Z(d[13]) );
  MUX2_X1 U766 ( .A(n1670), .B(n750), .S(n1546), .Z(n751) );
  MUX2_X1 U767 ( .A(n751), .B(n1663), .S(n1568), .Z(n752) );
  MUX2_X1 U768 ( .A(addr[0]), .B(n1671), .S(n1549), .Z(n753) );
  MUX2_X1 U769 ( .A(n577), .B(n1849), .S(n1520), .Z(n754) );
  MUX2_X1 U770 ( .A(n754), .B(n632), .S(n1550), .Z(n755) );
  MUX2_X1 U771 ( .A(n755), .B(n753), .S(n1568), .Z(n756) );
  MUX2_X1 U772 ( .A(n756), .B(n752), .S(n458), .Z(n757) );
  MUX2_X1 U774 ( .A(n757), .B(n758), .S(n1578), .Z(d[14]) );
  MUX2_X1 U776 ( .A(n760), .B(n1838), .S(n1520), .Z(n761) );
  MUX2_X1 U777 ( .A(n443), .B(n1813), .S(n1520), .Z(n762) );
  MUX2_X1 U778 ( .A(n762), .B(n761), .S(n458), .Z(n763) );
  MUX2_X1 U780 ( .A(n763), .B(n764), .S(n1552), .Z(n766) );
  MUX2_X1 U781 ( .A(n1744), .B(n1791), .S(n1520), .Z(n767) );
  MUX2_X1 U782 ( .A(n1761), .B(n1777), .S(n1520), .Z(n768) );
  MUX2_X1 U783 ( .A(n768), .B(n767), .S(n461), .Z(n769) );
  MUX2_X1 U784 ( .A(n1756), .B(n573), .S(n1520), .Z(n770) );
  MUX2_X1 U785 ( .A(n1797), .B(n539), .S(n1520), .Z(n771) );
  MUX2_X1 U786 ( .A(n771), .B(n770), .S(n458), .Z(n772) );
  MUX2_X1 U787 ( .A(n772), .B(n769), .S(n1551), .Z(n773) );
  MUX2_X1 U788 ( .A(n773), .B(n766), .S(n1568), .Z(n774) );
  MUX2_X1 U789 ( .A(n1756), .B(n1805), .S(n1520), .Z(n775) );
  MUX2_X1 U791 ( .A(n1810), .B(n776), .S(n1520), .Z(n777) );
  MUX2_X1 U792 ( .A(n777), .B(n775), .S(n458), .Z(n778) );
  MUX2_X1 U793 ( .A(n1756), .B(n1839), .S(n1520), .Z(n779) );
  MUX2_X1 U794 ( .A(n1743), .B(n627), .S(n1520), .Z(n780) );
  MUX2_X1 U795 ( .A(n780), .B(n779), .S(n458), .Z(n781) );
  MUX2_X1 U796 ( .A(n781), .B(n778), .S(n1552), .Z(n782) );
  MUX2_X1 U797 ( .A(n1742), .B(n1762), .S(n1521), .Z(n783) );
  MUX2_X1 U798 ( .A(n1741), .B(n541), .S(n1521), .Z(n784) );
  MUX2_X1 U799 ( .A(n784), .B(n783), .S(n458), .Z(n785) );
  MUX2_X1 U800 ( .A(n1786), .B(n540), .S(n1521), .Z(n786) );
  MUX2_X1 U801 ( .A(n569), .B(n1838), .S(n1521), .Z(n787) );
  MUX2_X1 U802 ( .A(n787), .B(n786), .S(n458), .Z(n788) );
  MUX2_X1 U803 ( .A(n788), .B(n785), .S(n1547), .Z(n789) );
  MUX2_X1 U804 ( .A(n789), .B(n782), .S(n1568), .Z(n790) );
  MUX2_X1 U805 ( .A(n790), .B(n774), .S(n1578), .Z(d[17]) );
  MUX2_X1 U806 ( .A(n597), .B(n1564), .S(n1521), .Z(n791) );
  MUX2_X1 U807 ( .A(n1834), .B(n539), .S(n1521), .Z(n792) );
  MUX2_X1 U808 ( .A(n1811), .B(n555), .S(addr[6]), .Z(n793) );
  MUX2_X1 U810 ( .A(n793), .B(n794), .S(n1521), .Z(n795) );
  MUX2_X1 U812 ( .A(n795), .B(n796), .S(n459), .Z(n797) );
  MUX2_X1 U813 ( .A(n1795), .B(n1807), .S(n1567), .Z(n798) );
  MUX2_X1 U814 ( .A(n1797), .B(n1760), .S(addr[6]), .Z(n799) );
  MUX2_X1 U815 ( .A(n799), .B(n798), .S(n1521), .Z(n800) );
  MUX2_X1 U816 ( .A(n1824), .B(n1774), .S(n1567), .Z(n801) );
  MUX2_X1 U817 ( .A(n586), .B(n1804), .S(addr[6]), .Z(n802) );
  MUX2_X1 U818 ( .A(n802), .B(n801), .S(n1521), .Z(n803) );
  MUX2_X1 U819 ( .A(n803), .B(n800), .S(n459), .Z(n804) );
  MUX2_X1 U820 ( .A(n804), .B(n797), .S(n1547), .Z(n805) );
  MUX2_X1 U821 ( .A(n532), .B(n572), .S(addr[6]), .Z(n806) );
  MUX2_X1 U823 ( .A(n806), .B(n807), .S(n1521), .Z(n808) );
  MUX2_X1 U824 ( .A(n531), .B(n1788), .S(addr[6]), .Z(n809) );
  MUX2_X1 U825 ( .A(n1743), .B(n1842), .S(addr[6]), .Z(n810) );
  MUX2_X1 U826 ( .A(n810), .B(n809), .S(n1521), .Z(n811) );
  MUX2_X1 U827 ( .A(n811), .B(n808), .S(n459), .Z(n812) );
  MUX2_X1 U828 ( .A(n589), .B(n1794), .S(addr[6]), .Z(n813) );
  MUX2_X1 U829 ( .A(n1838), .B(n1760), .S(addr[6]), .Z(n814) );
  MUX2_X1 U830 ( .A(n814), .B(n813), .S(n1521), .Z(n815) );
  MUX2_X1 U832 ( .A(n1756), .B(n816), .S(n1521), .Z(n818) );
  MUX2_X1 U833 ( .A(n818), .B(n815), .S(n459), .Z(n819) );
  MUX2_X1 U834 ( .A(n819), .B(n812), .S(n1546), .Z(n820) );
  MUX2_X1 U835 ( .A(n820), .B(n805), .S(n1578), .Z(d[18]) );
  MUX2_X1 U836 ( .A(n601), .B(n629), .S(n1564), .Z(n821) );
  MUX2_X1 U837 ( .A(n1772), .B(n1781), .S(addr[6]), .Z(n822) );
  MUX2_X1 U839 ( .A(n822), .B(n823), .S(n1521), .Z(n824) );
  MUX2_X1 U841 ( .A(n824), .B(n825), .S(n459), .Z(n826) );
  MUX2_X1 U842 ( .A(n1808), .B(n1776), .S(addr[6]), .Z(n827) );
  MUX2_X1 U843 ( .A(n1817), .B(n531), .S(addr[6]), .Z(n828) );
  MUX2_X1 U844 ( .A(n828), .B(n827), .S(n1521), .Z(n829) );
  MUX2_X1 U845 ( .A(n1850), .B(n1814), .S(addr[6]), .Z(n830) );
  MUX2_X1 U846 ( .A(n1754), .B(n1834), .S(addr[6]), .Z(n831) );
  MUX2_X1 U847 ( .A(n831), .B(n830), .S(n1521), .Z(n832) );
  MUX2_X1 U848 ( .A(n832), .B(n829), .S(n459), .Z(n833) );
  MUX2_X1 U849 ( .A(n833), .B(n826), .S(n1552), .Z(n834) );
  MUX2_X1 U850 ( .A(n1793), .B(n1786), .S(n1567), .Z(n835) );
  MUX2_X1 U852 ( .A(n835), .B(n836), .S(n1521), .Z(n838) );
  MUX2_X1 U853 ( .A(addr[2]), .B(n1854), .S(addr[6]), .Z(n839) );
  MUX2_X1 U854 ( .A(n1786), .B(n573), .S(n1567), .Z(n840) );
  MUX2_X1 U855 ( .A(n840), .B(n839), .S(n1521), .Z(n841) );
  MUX2_X1 U856 ( .A(n841), .B(n838), .S(n459), .Z(n842) );
  MUX2_X1 U857 ( .A(n1801), .B(n1817), .S(n1567), .Z(n843) );
  MUX2_X1 U859 ( .A(n843), .B(n844), .S(n1522), .Z(n845) );
  MUX2_X1 U860 ( .A(n529), .B(n1776), .S(n1567), .Z(n846) );
  MUX2_X1 U861 ( .A(n1764), .B(n1821), .S(n1567), .Z(n847) );
  MUX2_X1 U862 ( .A(n847), .B(n846), .S(n1522), .Z(n848) );
  MUX2_X1 U863 ( .A(n848), .B(n845), .S(n459), .Z(n849) );
  MUX2_X1 U864 ( .A(n849), .B(n842), .S(n1552), .Z(n850) );
  MUX2_X1 U865 ( .A(n850), .B(n834), .S(n1578), .Z(d[19]) );
  MUX2_X1 U866 ( .A(n1674), .B(n1792), .S(n1522), .Z(n851) );
  MUX2_X1 U867 ( .A(n1750), .B(n1764), .S(n1522), .Z(n852) );
  MUX2_X1 U868 ( .A(n852), .B(n851), .S(n459), .Z(n853) );
  MUX2_X1 U870 ( .A(n853), .B(n854), .S(n1552), .Z(n856) );
  MUX2_X1 U871 ( .A(n1779), .B(n760), .S(n1522), .Z(n857) );
  MUX2_X1 U872 ( .A(n435), .B(n410), .S(n1522), .Z(n858) );
  MUX2_X1 U873 ( .A(n858), .B(n857), .S(n459), .Z(n859) );
  MUX2_X1 U874 ( .A(n1778), .B(n1807), .S(n1522), .Z(n860) );
  MUX2_X1 U875 ( .A(n575), .B(n557), .S(n1522), .Z(n861) );
  MUX2_X1 U876 ( .A(n861), .B(n860), .S(n459), .Z(n862) );
  MUX2_X1 U877 ( .A(n862), .B(n859), .S(n1552), .Z(n863) );
  MUX2_X1 U878 ( .A(n863), .B(n856), .S(n1567), .Z(n864) );
  MUX2_X1 U879 ( .A(n1843), .B(n581), .S(n1522), .Z(n865) );
  MUX2_X1 U880 ( .A(n1759), .B(n1802), .S(n1522), .Z(n866) );
  MUX2_X1 U881 ( .A(n866), .B(n865), .S(n459), .Z(n867) );
  MUX2_X1 U882 ( .A(n525), .B(n1853), .S(n1522), .Z(n868) );
  MUX2_X1 U884 ( .A(n869), .B(n868), .S(n459), .Z(n870) );
  MUX2_X1 U885 ( .A(n870), .B(n867), .S(n1552), .Z(n871) );
  MUX2_X1 U886 ( .A(n547), .B(n1759), .S(n1522), .Z(n872) );
  MUX2_X1 U888 ( .A(n872), .B(n873), .S(n459), .Z(n874) );
  MUX2_X1 U889 ( .A(n1761), .B(n1767), .S(n1522), .Z(n875) );
  MUX2_X1 U890 ( .A(n1815), .B(n1674), .S(n1522), .Z(n876) );
  MUX2_X1 U891 ( .A(n876), .B(n875), .S(n459), .Z(n877) );
  MUX2_X1 U892 ( .A(n877), .B(n874), .S(n1552), .Z(n878) );
  MUX2_X1 U893 ( .A(n878), .B(n871), .S(n1567), .Z(n879) );
  MUX2_X1 U894 ( .A(n879), .B(n864), .S(n1578), .Z(d[1]) );
  MUX2_X1 U895 ( .A(n527), .B(n538), .S(n459), .Z(n880) );
  MUX2_X1 U896 ( .A(n526), .B(n520), .S(n459), .Z(n881) );
  MUX2_X1 U897 ( .A(n881), .B(n880), .S(n1522), .Z(n882) );
  MUX2_X1 U899 ( .A(n882), .B(n883), .S(n1543), .Z(n885) );
  MUX2_X1 U900 ( .A(n1741), .B(n1831), .S(n459), .Z(n886) );
  MUX2_X1 U901 ( .A(n563), .B(n542), .S(n460), .Z(n887) );
  MUX2_X1 U902 ( .A(n887), .B(n886), .S(n1522), .Z(n888) );
  MUX2_X1 U903 ( .A(n1820), .B(n523), .S(n460), .Z(n889) );
  MUX2_X1 U904 ( .A(n443), .B(n889), .S(n1522), .Z(n890) );
  MUX2_X1 U905 ( .A(n890), .B(n888), .S(n1552), .Z(n891) );
  MUX2_X1 U906 ( .A(n891), .B(n885), .S(n1567), .Z(n892) );
  MUX2_X1 U907 ( .A(n1789), .B(n1784), .S(n460), .Z(n893) );
  MUX2_X1 U908 ( .A(n1782), .B(n603), .S(n460), .Z(n894) );
  MUX2_X1 U909 ( .A(n894), .B(n893), .S(n1522), .Z(n895) );
  MUX2_X1 U910 ( .A(n562), .B(n591), .S(n460), .Z(n896) );
  MUX2_X1 U912 ( .A(n517), .B(n897), .S(n460), .Z(n898) );
  MUX2_X1 U913 ( .A(n898), .B(n896), .S(n1523), .Z(n899) );
  MUX2_X1 U914 ( .A(n899), .B(n895), .S(n1552), .Z(n900) );
  MUX2_X1 U915 ( .A(n557), .B(n502), .S(n460), .Z(n901) );
  MUX2_X1 U916 ( .A(n901), .B(n555), .S(n1523), .Z(n902) );
  MUX2_X1 U917 ( .A(n1785), .B(n1745), .S(n460), .Z(n903) );
  MUX2_X1 U918 ( .A(n1775), .B(n556), .S(n460), .Z(n904) );
  MUX2_X1 U919 ( .A(n904), .B(n903), .S(n1523), .Z(n905) );
  MUX2_X1 U920 ( .A(n905), .B(n902), .S(n1552), .Z(n906) );
  MUX2_X1 U921 ( .A(n906), .B(n900), .S(n1567), .Z(n907) );
  MUX2_X1 U922 ( .A(n907), .B(n892), .S(n1578), .Z(d[20]) );
  MUX2_X1 U923 ( .A(n1798), .B(n523), .S(n460), .Z(n908) );
  MUX2_X1 U924 ( .A(n1779), .B(n608), .S(n460), .Z(n909) );
  MUX2_X1 U926 ( .A(n910), .B(n909), .S(n1523), .Z(n911) );
  MUX2_X1 U928 ( .A(n911), .B(n912), .S(n1551), .Z(n913) );
  MUX2_X1 U929 ( .A(n1843), .B(n548), .S(n460), .Z(n914) );
  MUX2_X1 U930 ( .A(n1853), .B(n1767), .S(n460), .Z(n915) );
  MUX2_X1 U931 ( .A(n915), .B(n914), .S(n1523), .Z(n916) );
  MUX2_X1 U932 ( .A(n1796), .B(n1815), .S(n460), .Z(n917) );
  MUX2_X1 U933 ( .A(n563), .B(n760), .S(n460), .Z(n918) );
  MUX2_X1 U934 ( .A(n918), .B(n917), .S(n1523), .Z(n919) );
  MUX2_X1 U935 ( .A(n919), .B(n916), .S(n1546), .Z(n920) );
  MUX2_X1 U936 ( .A(n920), .B(n913), .S(n1567), .Z(n921) );
  MUX2_X1 U937 ( .A(n548), .B(n1818), .S(n460), .Z(n922) );
  MUX2_X1 U938 ( .A(n554), .B(n1793), .S(n460), .Z(n923) );
  MUX2_X1 U939 ( .A(n923), .B(n922), .S(n1523), .Z(n924) );
  MUX2_X1 U940 ( .A(n1803), .B(n593), .S(n460), .Z(n925) );
  MUX2_X1 U941 ( .A(n410), .B(n517), .S(n461), .Z(n926) );
  MUX2_X1 U942 ( .A(n926), .B(n925), .S(n1523), .Z(n927) );
  MUX2_X1 U943 ( .A(n927), .B(n924), .S(n1545), .Z(n928) );
  MUX2_X1 U944 ( .A(n1760), .B(n583), .S(n461), .Z(n929) );
  MUX2_X1 U945 ( .A(n929), .B(n1806), .S(n1523), .Z(n930) );
  MUX2_X1 U946 ( .A(n562), .B(n550), .S(n461), .Z(n931) );
  MUX2_X1 U948 ( .A(n932), .B(n931), .S(n1523), .Z(n933) );
  MUX2_X1 U949 ( .A(n933), .B(n930), .S(n1545), .Z(n934) );
  MUX2_X1 U950 ( .A(n934), .B(n928), .S(n1567), .Z(n935) );
  MUX2_X1 U951 ( .A(n935), .B(n921), .S(n1578), .Z(d[21]) );
  MUX2_X1 U952 ( .A(n602), .B(n1800), .S(n461), .Z(n936) );
  MUX2_X1 U953 ( .A(n583), .B(n1787), .S(n1523), .Z(n937) );
  MUX2_X1 U954 ( .A(n555), .B(n601), .S(n1523), .Z(n938) );
  MUX2_X1 U955 ( .A(n938), .B(n937), .S(n461), .Z(n939) );
  MUX2_X1 U957 ( .A(n939), .B(n940), .S(n1545), .Z(n941) );
  MUX2_X1 U958 ( .A(n1808), .B(n542), .S(n1523), .Z(n942) );
  MUX2_X1 U959 ( .A(n608), .B(n573), .S(n1523), .Z(n943) );
  MUX2_X1 U960 ( .A(n943), .B(n942), .S(n461), .Z(n944) );
  MUX2_X1 U961 ( .A(n776), .B(n564), .S(n1523), .Z(n945) );
  MUX2_X1 U962 ( .A(n570), .B(n1834), .S(n1523), .Z(n946) );
  MUX2_X1 U963 ( .A(n946), .B(n945), .S(n461), .Z(n947) );
  MUX2_X1 U964 ( .A(n947), .B(n944), .S(n1545), .Z(n948) );
  MUX2_X1 U965 ( .A(n948), .B(n941), .S(n1567), .Z(n949) );
  MUX2_X1 U966 ( .A(n527), .B(n588), .S(n1523), .Z(n950) );
  MUX2_X1 U967 ( .A(n1825), .B(n1762), .S(n1523), .Z(n951) );
  MUX2_X1 U968 ( .A(n951), .B(n950), .S(n461), .Z(n952) );
  MUX2_X1 U969 ( .A(n1829), .B(n565), .S(n1524), .Z(n953) );
  MUX2_X1 U970 ( .A(n1845), .B(n1759), .S(n1524), .Z(n954) );
  MUX2_X1 U971 ( .A(n954), .B(n953), .S(n461), .Z(n955) );
  MUX2_X1 U972 ( .A(n955), .B(n952), .S(n1545), .Z(n956) );
  MUX2_X1 U973 ( .A(n1802), .B(n595), .S(n1524), .Z(n957) );
  MUX2_X1 U974 ( .A(n1799), .B(n1790), .S(n1524), .Z(n958) );
  MUX2_X1 U975 ( .A(n958), .B(n957), .S(n461), .Z(n959) );
  MUX2_X1 U976 ( .A(n522), .B(n1743), .S(n1524), .Z(n960) );
  MUX2_X1 U977 ( .A(n526), .B(n445), .S(n1524), .Z(n961) );
  MUX2_X1 U978 ( .A(n961), .B(n960), .S(n461), .Z(n962) );
  MUX2_X1 U979 ( .A(n962), .B(n959), .S(n1545), .Z(n963) );
  MUX2_X1 U980 ( .A(n963), .B(n956), .S(n1567), .Z(n964) );
  MUX2_X1 U981 ( .A(n964), .B(n949), .S(n1578), .Z(d[22]) );
  MUX2_X1 U982 ( .A(n1812), .B(addr[2]), .S(n461), .Z(n965) );
  MUX2_X1 U983 ( .A(n591), .B(n1754), .S(n1524), .Z(n966) );
  MUX2_X1 U985 ( .A(n967), .B(n966), .S(n461), .Z(n968) );
  MUX2_X1 U987 ( .A(n968), .B(n969), .S(n1545), .Z(n970) );
  MUX2_X1 U988 ( .A(n1821), .B(n520), .S(n1524), .Z(n971) );
  MUX2_X1 U989 ( .A(n530), .B(n1797), .S(n1524), .Z(n972) );
  MUX2_X1 U990 ( .A(n972), .B(n971), .S(n461), .Z(n973) );
  MUX2_X1 U991 ( .A(n544), .B(n1754), .S(n461), .Z(n974) );
  MUX2_X1 U992 ( .A(n547), .B(n974), .S(n428), .Z(n975) );
  MUX2_X1 U993 ( .A(n975), .B(n973), .S(n1545), .Z(n976) );
  MUX2_X1 U994 ( .A(n976), .B(n970), .S(n1567), .Z(n977) );
  MUX2_X1 U995 ( .A(n1783), .B(n602), .S(n1524), .Z(n978) );
  MUX2_X1 U996 ( .A(n1780), .B(n565), .S(n1524), .Z(n979) );
  MUX2_X1 U997 ( .A(n979), .B(n978), .S(n461), .Z(n980) );
  MUX2_X1 U998 ( .A(n571), .B(n583), .S(n1524), .Z(n981) );
  MUX2_X1 U999 ( .A(addr[2]), .B(n586), .S(n1524), .Z(n982) );
  MUX2_X1 U1000 ( .A(n982), .B(n981), .S(n461), .Z(n983) );
  MUX2_X1 U1001 ( .A(n983), .B(n980), .S(n1543), .Z(n984) );
  MUX2_X1 U1002 ( .A(n1830), .B(n606), .S(n1524), .Z(n985) );
  MUX2_X1 U1003 ( .A(n571), .B(n1775), .S(n1524), .Z(n986) );
  MUX2_X1 U1004 ( .A(n986), .B(n985), .S(n453), .Z(n987) );
  MUX2_X1 U1005 ( .A(n1777), .B(n612), .S(n1524), .Z(n988) );
  MUX2_X1 U1006 ( .A(n1830), .B(n572), .S(n1524), .Z(n989) );
  MUX2_X1 U1007 ( .A(n989), .B(n988), .S(n460), .Z(n990) );
  MUX2_X1 U1008 ( .A(n990), .B(n987), .S(n1545), .Z(n991) );
  MUX2_X1 U1009 ( .A(n991), .B(n984), .S(n1567), .Z(n992) );
  MUX2_X1 U1010 ( .A(n992), .B(n977), .S(n1578), .Z(d[23]) );
  MUX2_X1 U1013 ( .A(n994), .B(n993), .S(n1524), .Z(n995) );
  MUX2_X1 U1014 ( .A(n1755), .B(n615), .S(n1578), .Z(n996) );
  MUX2_X1 U1016 ( .A(n996), .B(n997), .S(n504), .Z(n998) );
  MUX2_X1 U1017 ( .A(n998), .B(n995), .S(n459), .Z(n999) );
  MUX2_X1 U1018 ( .A(n579), .B(n609), .S(n1577), .Z(n1000) );
  MUX2_X1 U1019 ( .A(n1840), .B(n1745), .S(n1578), .Z(n1001) );
  MUX2_X1 U1020 ( .A(n1001), .B(n1000), .S(n504), .Z(n1002) );
  MUX2_X1 U1021 ( .A(n566), .B(n629), .S(n1577), .Z(n1003) );
  MUX2_X1 U1022 ( .A(n1756), .B(n584), .S(n1577), .Z(n1004) );
  MUX2_X1 U1023 ( .A(n1004), .B(n1003), .S(n504), .Z(n1005) );
  MUX2_X1 U1024 ( .A(n1005), .B(n1002), .S(n455), .Z(n1006) );
  MUX2_X1 U1025 ( .A(n1006), .B(n999), .S(n1545), .Z(n1007) );
  MUX2_X1 U1026 ( .A(n537), .B(n4870), .S(n1577), .Z(n1008) );
  MUX2_X1 U1027 ( .A(n593), .B(n617), .S(n1577), .Z(n1009) );
  MUX2_X1 U1028 ( .A(n1009), .B(n1008), .S(n504), .Z(n1010) );
  MUX2_X1 U1029 ( .A(n1813), .B(n562), .S(n1577), .Z(n1011) );
  MUX2_X1 U1030 ( .A(n1752), .B(n1747), .S(n1577), .Z(n1012) );
  MUX2_X1 U1031 ( .A(n1012), .B(n1011), .S(n504), .Z(n1013) );
  MUX2_X1 U1032 ( .A(n1013), .B(n1010), .S(n462), .Z(n1014) );
  MUX2_X1 U1033 ( .A(n564), .B(n1746), .S(n1577), .Z(n1015) );
  MUX2_X1 U1034 ( .A(n897), .B(n1769), .S(n1577), .Z(n1016) );
  MUX2_X1 U1035 ( .A(n1016), .B(n1015), .S(n505), .Z(n1017) );
  MUX2_X1 U1036 ( .A(n615), .B(n1768), .S(n1577), .Z(n1018) );
  MUX2_X1 U1037 ( .A(n555), .B(addr[0]), .S(n1577), .Z(n1019) );
  MUX2_X1 U1038 ( .A(n1019), .B(n1018), .S(n504), .Z(n1020) );
  MUX2_X1 U1039 ( .A(n1020), .B(n1017), .S(n457), .Z(n1021) );
  MUX2_X1 U1040 ( .A(n1021), .B(n1014), .S(n1545), .Z(n1022) );
  MUX2_X1 U1041 ( .A(n1022), .B(n1007), .S(n1567), .Z(d[24]) );
  MUX2_X1 U1042 ( .A(n601), .B(n1826), .S(n505), .Z(n1023) );
  MUX2_X1 U1044 ( .A(n1024), .B(n1023), .S(n456), .Z(n1025) );
  MUX2_X1 U1046 ( .A(n1025), .B(n1026), .S(n1552), .Z(n1028) );
  MUX2_X1 U1047 ( .A(n557), .B(n533), .S(n510), .Z(n1029) );
  MUX2_X1 U1048 ( .A(n561), .B(n1789), .S(n510), .Z(n1030) );
  MUX2_X1 U1049 ( .A(n1030), .B(n1029), .S(n456), .Z(n1031) );
  MUX2_X1 U1050 ( .A(n1839), .B(n573), .S(n510), .Z(n1032) );
  MUX2_X1 U1051 ( .A(n1672), .B(n1032), .S(n458), .Z(n1033) );
  MUX2_X1 U1052 ( .A(n1033), .B(n1031), .S(n1545), .Z(n1034) );
  MUX2_X1 U1053 ( .A(n1034), .B(n1028), .S(n1566), .Z(n1035) );
  MUX2_X1 U1054 ( .A(n613), .B(n576), .S(n510), .Z(n1036) );
  MUX2_X1 U1055 ( .A(n605), .B(n1841), .S(n510), .Z(n1037) );
  MUX2_X1 U1056 ( .A(n1037), .B(n1036), .S(n462), .Z(n1038) );
  MUX2_X1 U1057 ( .A(n1820), .B(n1824), .S(n510), .Z(n1039) );
  MUX2_X1 U1058 ( .A(n1818), .B(n1795), .S(n510), .Z(n1040) );
  MUX2_X1 U1059 ( .A(n1040), .B(n1039), .S(n454), .Z(n1041) );
  MUX2_X1 U1060 ( .A(n1041), .B(n1038), .S(n1552), .Z(n1042) );
  MUX2_X1 U1061 ( .A(n1805), .B(n598), .S(n510), .Z(n1043) );
  MUX2_X1 U1062 ( .A(n1826), .B(n566), .S(n510), .Z(n1044) );
  MUX2_X1 U1063 ( .A(n1044), .B(n1043), .S(n461), .Z(n1045) );
  MUX2_X1 U1064 ( .A(n592), .B(n897), .S(n510), .Z(n1046) );
  MUX2_X1 U1065 ( .A(n535), .B(n567), .S(n510), .Z(n1047) );
  MUX2_X1 U1066 ( .A(n1047), .B(n1046), .S(n451), .Z(n1048) );
  MUX2_X1 U1067 ( .A(n1048), .B(n1045), .S(n1545), .Z(n1049) );
  MUX2_X1 U1068 ( .A(n1049), .B(n1042), .S(n1567), .Z(n1050) );
  MUX2_X1 U1069 ( .A(n1050), .B(n1035), .S(n1577), .Z(d[25]) );
  MUX2_X1 U1070 ( .A(n536), .B(n628), .S(n456), .Z(n1051) );
  MUX2_X1 U1071 ( .A(n612), .B(n1833), .S(n510), .Z(n1052) );
  MUX2_X1 U1072 ( .A(n493), .B(n601), .S(n5090), .Z(n1053) );
  MUX2_X1 U1073 ( .A(n1053), .B(n1052), .S(n456), .Z(n1054) );
  MUX2_X1 U1075 ( .A(n1054), .B(n1055), .S(n1546), .Z(n1056) );
  MUX2_X1 U1076 ( .A(n1809), .B(n1802), .S(n5090), .Z(n1057) );
  MUX2_X1 U1077 ( .A(n566), .B(n1827), .S(n5090), .Z(n1058) );
  MUX2_X1 U1078 ( .A(n1058), .B(n1057), .S(n456), .Z(n1059) );
  MUX2_X1 U1079 ( .A(n1776), .B(n567), .S(n5090), .Z(n1060) );
  MUX2_X1 U1081 ( .A(n1061), .B(n1060), .S(n462), .Z(n1062) );
  MUX2_X1 U1082 ( .A(n1062), .B(n1059), .S(n1545), .Z(n1063) );
  MUX2_X1 U1083 ( .A(n1063), .B(n1056), .S(n1566), .Z(n1064) );
  MUX2_X1 U1084 ( .A(n1748), .B(n619), .S(n5090), .Z(n1065) );
  MUX2_X1 U1085 ( .A(n1846), .B(n523), .S(n5090), .Z(n1066) );
  MUX2_X1 U1086 ( .A(n1066), .B(n1065), .S(n456), .Z(n1067) );
  MUX2_X1 U1087 ( .A(n602), .B(n629), .S(n5090), .Z(n1068) );
  MUX2_X1 U1088 ( .A(n1068), .B(n1070), .S(n462), .Z(n1069) );
  MUX2_X1 U1089 ( .A(n1069), .B(n1067), .S(n1545), .Z(n1071) );
  MUX2_X1 U1090 ( .A(n1742), .B(n1779), .S(n5090), .Z(n1072) );
  MUX2_X1 U1091 ( .A(n596), .B(n560), .S(n5090), .Z(n1073) );
  MUX2_X1 U1092 ( .A(n1073), .B(n1072), .S(n462), .Z(n1074) );
  MUX2_X1 U1093 ( .A(n599), .B(n1820), .S(n5090), .Z(n1075) );
  MUX2_X1 U1094 ( .A(n1771), .B(n523), .S(n5090), .Z(n1076) );
  MUX2_X1 U1095 ( .A(n1076), .B(n1075), .S(n462), .Z(n1077) );
  MUX2_X1 U1096 ( .A(n1077), .B(n1074), .S(n1545), .Z(n1078) );
  MUX2_X1 U1097 ( .A(n1078), .B(n1071), .S(n1567), .Z(n1079) );
  MUX2_X1 U1098 ( .A(n1079), .B(n1064), .S(n1577), .Z(d[26]) );
  MUX2_X1 U1099 ( .A(n593), .B(n581), .S(n5090), .Z(n1080) );
  MUX2_X1 U1100 ( .A(addr[0]), .B(n612), .S(n5090), .Z(n1081) );
  MUX2_X1 U1101 ( .A(n1081), .B(n1080), .S(n462), .Z(n1082) );
  MUX2_X1 U1103 ( .A(n1082), .B(n1083), .S(n1547), .Z(n1085) );
  MUX2_X1 U1105 ( .A(n1809), .B(n1086), .S(n428), .Z(n1087) );
  MUX2_X1 U1106 ( .A(n1798), .B(n581), .S(n5090), .Z(n1088) );
  MUX2_X1 U1107 ( .A(n1808), .B(n536), .S(n5090), .Z(n1089) );
  MUX2_X1 U1108 ( .A(n1089), .B(n1088), .S(n462), .Z(n1090) );
  MUX2_X1 U1109 ( .A(n1090), .B(n1087), .S(n1547), .Z(n1091) );
  MUX2_X1 U1110 ( .A(n1091), .B(n1085), .S(n1566), .Z(n1092) );
  MUX2_X1 U1111 ( .A(n410), .B(n1826), .S(n5090), .Z(n1093) );
  MUX2_X1 U1113 ( .A(n1093), .B(n1094), .S(n462), .Z(n1095) );
  MUX2_X1 U1114 ( .A(n410), .B(n1805), .S(n5090), .Z(n1096) );
  MUX2_X1 U1115 ( .A(n598), .B(n557), .S(n5090), .Z(n1097) );
  MUX2_X1 U1116 ( .A(n1097), .B(n1096), .S(n462), .Z(n1098) );
  MUX2_X1 U1117 ( .A(n1098), .B(n1095), .S(n1552), .Z(n1099) );
  MUX2_X1 U1118 ( .A(n1841), .B(n1759), .S(n508), .Z(n1100) );
  MUX2_X1 U1119 ( .A(n548), .B(n620), .S(n508), .Z(n1101) );
  MUX2_X1 U1120 ( .A(n1101), .B(n1100), .S(n462), .Z(n1102) );
  MUX2_X1 U1121 ( .A(n565), .B(n545), .S(n508), .Z(n1103) );
  MUX2_X1 U1122 ( .A(n1749), .B(n1825), .S(n508), .Z(n1104) );
  MUX2_X1 U1123 ( .A(n1104), .B(n1103), .S(n462), .Z(n1105) );
  MUX2_X1 U1124 ( .A(n1105), .B(n1102), .S(n1552), .Z(n1106) );
  MUX2_X1 U1125 ( .A(n1106), .B(n1099), .S(n1566), .Z(n1107) );
  MUX2_X1 U1126 ( .A(n1107), .B(n1092), .S(n1577), .Z(d[27]) );
  MUX2_X1 U1127 ( .A(n479), .B(n624), .S(n1546), .Z(n1108) );
  MUX2_X1 U1128 ( .A(n623), .B(n1821), .S(n1547), .Z(n1109) );
  MUX2_X1 U1130 ( .A(n1110), .B(addr[0]), .S(n462), .Z(n1111) );
  MUX2_X1 U1132 ( .A(n1112), .B(n623), .S(n462), .Z(n1113) );
  MUX2_X1 U1133 ( .A(n1113), .B(n1111), .S(n1552), .Z(n1114) );
  MUX2_X1 U1135 ( .A(n1114), .B(n1115), .S(n1566), .Z(n1117) );
  MUX2_X1 U1136 ( .A(n539), .B(n1826), .S(n508), .Z(n1118) );
  MUX2_X1 U1137 ( .A(n1118), .B(n1667), .S(n462), .Z(n1119) );
  MUX2_X1 U1138 ( .A(n1809), .B(n567), .S(n508), .Z(n1120) );
  MUX2_X1 U1139 ( .A(n551), .B(n1794), .S(n508), .Z(n1121) );
  MUX2_X1 U1140 ( .A(n1121), .B(n1120), .S(n462), .Z(n1122) );
  MUX2_X1 U1141 ( .A(n1122), .B(n1119), .S(n1552), .Z(n1123) );
  MUX2_X1 U1142 ( .A(n523), .B(n567), .S(n508), .Z(n1124) );
  MUX2_X1 U1143 ( .A(n590), .B(n1789), .S(n508), .Z(n1125) );
  MUX2_X1 U1144 ( .A(n1125), .B(n1124), .S(n462), .Z(n1126) );
  MUX2_X1 U1145 ( .A(n533), .B(n606), .S(n508), .Z(n1127) );
  MUX2_X1 U1146 ( .A(n443), .B(n1768), .S(n508), .Z(n1128) );
  MUX2_X1 U1147 ( .A(n1128), .B(n1127), .S(n462), .Z(n1129) );
  MUX2_X1 U1148 ( .A(n1129), .B(n1126), .S(n1551), .Z(n1130) );
  MUX2_X1 U1149 ( .A(n1130), .B(n1123), .S(n1566), .Z(n1131) );
  MUX2_X1 U1150 ( .A(n1131), .B(n1117), .S(n1578), .Z(d[28]) );
  MUX2_X1 U1151 ( .A(n1585), .B(n431), .S(n462), .Z(n1132) );
  MUX2_X1 U1153 ( .A(n432), .B(n1133), .S(n463), .Z(n1134) );
  MUX2_X1 U1154 ( .A(n1134), .B(n1132), .S(n510), .Z(n1135) );
  MUX2_X1 U1155 ( .A(n536), .B(n1820), .S(n1577), .Z(n1136) );
  MUX2_X1 U1157 ( .A(n1136), .B(n1137), .S(n462), .Z(n1138) );
  MUX2_X1 U1159 ( .A(n1139), .B(n1138), .S(n508), .Z(n1140) );
  MUX2_X1 U1160 ( .A(n1140), .B(n1135), .S(n1544), .Z(n1141) );
  MUX2_X1 U1161 ( .A(n1832), .B(n1834), .S(n1577), .Z(n1142) );
  MUX2_X1 U1163 ( .A(n1142), .B(n1143), .S(n463), .Z(n1144) );
  MUX2_X1 U1164 ( .A(n1798), .B(n445), .S(n1576), .Z(n1145) );
  MUX2_X1 U1165 ( .A(n1145), .B(n546), .S(n463), .Z(n1146) );
  MUX2_X1 U1166 ( .A(n1146), .B(n1144), .S(n508), .Z(n1147) );
  MUX2_X1 U1167 ( .A(n1819), .B(n551), .S(n1577), .Z(n1148) );
  MUX2_X1 U1168 ( .A(n594), .B(n446), .S(n1576), .Z(n1149) );
  MUX2_X1 U1169 ( .A(n1149), .B(n1148), .S(n463), .Z(n1150) );
  MUX2_X1 U1170 ( .A(n1854), .B(addr[0]), .S(n1577), .Z(n1151) );
  MUX2_X1 U1171 ( .A(n1812), .B(n445), .S(n1576), .Z(n1152) );
  MUX2_X1 U1172 ( .A(n1152), .B(n1151), .S(n463), .Z(n1153) );
  MUX2_X1 U1173 ( .A(n1153), .B(n1150), .S(n508), .Z(n1154) );
  MUX2_X1 U1174 ( .A(n1154), .B(n1147), .S(n1550), .Z(n1155) );
  MUX2_X1 U1175 ( .A(n1155), .B(n1141), .S(n1566), .Z(d[29]) );
  MUX2_X1 U1176 ( .A(n625), .B(n1835), .S(n463), .Z(n1156) );
  MUX2_X1 U1177 ( .A(n552), .B(n1752), .S(n463), .Z(n1157) );
  MUX2_X1 U1178 ( .A(n1157), .B(n1156), .S(n507), .Z(n1158) );
  MUX2_X1 U1180 ( .A(n1158), .B(n1159), .S(n1544), .Z(n1161) );
  MUX2_X1 U1181 ( .A(n587), .B(n610), .S(n462), .Z(n1162) );
  MUX2_X1 U1182 ( .A(n616), .B(n551), .S(n454), .Z(n1163) );
  MUX2_X1 U1183 ( .A(n1163), .B(n1162), .S(n507), .Z(n1164) );
  MUX2_X1 U1184 ( .A(n1741), .B(n582), .S(n451), .Z(n1165) );
  MUX2_X1 U1186 ( .A(n1165), .B(n1166), .S(n507), .Z(n1167) );
  MUX2_X1 U1187 ( .A(n1167), .B(n1164), .S(n1546), .Z(n1168) );
  MUX2_X1 U1188 ( .A(n1168), .B(n1161), .S(n1566), .Z(n1169) );
  MUX2_X1 U1189 ( .A(n549), .B(n585), .S(n450), .Z(n1170) );
  MUX2_X1 U1191 ( .A(n1170), .B(n1171), .S(n508), .Z(n1172) );
  MUX2_X1 U1192 ( .A(n1758), .B(n1769), .S(n451), .Z(n1173) );
  MUX2_X1 U1193 ( .A(n604), .B(n583), .S(n450), .Z(n1174) );
  MUX2_X1 U1194 ( .A(n1174), .B(n1173), .S(n507), .Z(n1175) );
  MUX2_X1 U1195 ( .A(n1175), .B(n1172), .S(n1546), .Z(n1176) );
  MUX2_X1 U1196 ( .A(n4870), .B(n493), .S(n451), .Z(n1177) );
  MUX2_X1 U1197 ( .A(n1742), .B(n1749), .S(n451), .Z(n1178) );
  MUX2_X1 U1198 ( .A(n1178), .B(n1177), .S(n507), .Z(n1179) );
  MUX2_X1 U1199 ( .A(n606), .B(n1823), .S(n451), .Z(n1180) );
  MUX2_X1 U1200 ( .A(n1180), .B(n1806), .S(n507), .Z(n1181) );
  MUX2_X1 U1201 ( .A(n1181), .B(n1179), .S(n1551), .Z(n1182) );
  MUX2_X1 U1202 ( .A(n1182), .B(n1176), .S(n1566), .Z(n1183) );
  MUX2_X1 U1203 ( .A(n1183), .B(n1169), .S(n1576), .Z(d[2]) );
  MUX2_X1 U1204 ( .A(addr[0]), .B(n569), .S(n507), .Z(n1184) );
  MUX2_X1 U1205 ( .A(n1184), .B(n529), .S(n1566), .Z(n1185) );
  MUX2_X1 U1206 ( .A(n435), .B(n1185), .S(n1546), .Z(n1186) );
  MUX2_X1 U1208 ( .A(n463), .B(n1187), .S(n1566), .Z(n1188) );
  MUX2_X1 U1209 ( .A(n443), .B(n1820), .S(n507), .Z(n1189) );
  MUX2_X1 U1211 ( .A(n1189), .B(n1190), .S(n451), .Z(n1191) );
  MUX2_X1 U1213 ( .A(n1191), .B(n1192), .S(n1566), .Z(n1193) );
  MUX2_X1 U1214 ( .A(n1671), .B(n623), .S(n451), .Z(n1194) );
  MUX2_X1 U1215 ( .A(n776), .B(n1792), .S(n507), .Z(n1195) );
  MUX2_X1 U1216 ( .A(n615), .B(n565), .S(n508), .Z(n1196) );
  MUX2_X1 U1217 ( .A(n1196), .B(n1195), .S(n451), .Z(n1197) );
  MUX2_X1 U1218 ( .A(n1197), .B(n1194), .S(n1566), .Z(n1198) );
  MUX2_X1 U1219 ( .A(n1198), .B(n1193), .S(n1546), .Z(n1199) );
  MUX2_X1 U1221 ( .A(n1199), .B(n1200), .S(n1576), .Z(d[30]) );
  MUX2_X1 U1222 ( .A(n1791), .B(n1752), .S(n507), .Z(n1201) );
  MUX2_X1 U1223 ( .A(n1201), .B(n1813), .S(n451), .Z(n1202) );
  MUX2_X1 U1224 ( .A(n620), .B(n1763), .S(n451), .Z(n1203) );
  MUX2_X1 U1226 ( .A(n1204), .B(n1203), .S(n507), .Z(n1205) );
  MUX2_X1 U1227 ( .A(n1205), .B(n1202), .S(n1546), .Z(n1206) );
  MUX2_X1 U1229 ( .A(n554), .B(n543), .S(n451), .Z(n1207) );
  MUX2_X1 U1230 ( .A(n563), .B(n620), .S(n451), .Z(n1208) );
  MUX2_X1 U1231 ( .A(n1208), .B(n1207), .S(n506), .Z(n1209) );
  MUX2_X1 U1232 ( .A(n1828), .B(n1834), .S(n451), .Z(n1210) );
  MUX2_X1 U1233 ( .A(n610), .B(n615), .S(n451), .Z(n1211) );
  MUX2_X1 U1234 ( .A(n1211), .B(n1210), .S(n508), .Z(n1212) );
  MUX2_X1 U1235 ( .A(n1212), .B(n1209), .S(n1546), .Z(n1213) );
  MUX2_X1 U1236 ( .A(n1213), .B(n1206), .S(n1566), .Z(n1214) );
  MUX2_X1 U1237 ( .A(n1791), .B(n606), .S(n451), .Z(n1215) );
  MUX2_X1 U1238 ( .A(n1811), .B(n1788), .S(n451), .Z(n1216) );
  MUX2_X1 U1239 ( .A(n1216), .B(n1215), .S(n506), .Z(n1217) );
  MUX2_X1 U1240 ( .A(n625), .B(n1820), .S(n451), .Z(n1218) );
  MUX2_X1 U1241 ( .A(n1783), .B(n1803), .S(n451), .Z(n1219) );
  MUX2_X1 U1242 ( .A(n1219), .B(n1218), .S(n507), .Z(n1220) );
  MUX2_X1 U1243 ( .A(n1220), .B(n1217), .S(n1546), .Z(n1221) );
  MUX2_X1 U1244 ( .A(n528), .B(n570), .S(n452), .Z(n1222) );
  MUX2_X1 U1245 ( .A(n610), .B(n1772), .S(n452), .Z(n1223) );
  MUX2_X1 U1246 ( .A(n1223), .B(n1222), .S(n506), .Z(n1224) );
  MUX2_X1 U1247 ( .A(n1829), .B(n614), .S(n452), .Z(n1225) );
  MUX2_X1 U1248 ( .A(n1757), .B(n1225), .S(n507), .Z(n1226) );
  MUX2_X1 U1249 ( .A(n1226), .B(n1224), .S(n1546), .Z(n1227) );
  MUX2_X1 U1250 ( .A(n1227), .B(n1221), .S(n1566), .Z(n1228) );
  MUX2_X1 U1251 ( .A(n1228), .B(n1214), .S(n1576), .Z(d[35]) );
  MUX2_X1 U1254 ( .A(n1230), .B(n1229), .S(n507), .Z(n1231) );
  MUX2_X1 U1255 ( .A(n1826), .B(n610), .S(n452), .Z(n1232) );
  MUX2_X1 U1256 ( .A(n1824), .B(n1769), .S(n452), .Z(n1233) );
  MUX2_X1 U1257 ( .A(n1233), .B(n1232), .S(n506), .Z(n1234) );
  MUX2_X1 U1258 ( .A(n1234), .B(n1231), .S(n1546), .Z(n1235) );
  MUX2_X1 U1259 ( .A(n1814), .B(n1775), .S(n452), .Z(n1236) );
  MUX2_X1 U1260 ( .A(n1752), .B(n1797), .S(n452), .Z(n1237) );
  MUX2_X1 U1261 ( .A(n1237), .B(n1236), .S(n507), .Z(n1238) );
  MUX2_X1 U1262 ( .A(n609), .B(n536), .S(n452), .Z(n1239) );
  MUX2_X1 U1263 ( .A(n532), .B(n589), .S(n452), .Z(n1240) );
  MUX2_X1 U1264 ( .A(n1240), .B(n1239), .S(n506), .Z(n1241) );
  MUX2_X1 U1265 ( .A(n1241), .B(n1238), .S(n1546), .Z(n1242) );
  MUX2_X1 U1266 ( .A(n1242), .B(n1235), .S(n1566), .Z(n1243) );
  MUX2_X1 U1267 ( .A(n541), .B(n577), .S(n452), .Z(n1244) );
  MUX2_X1 U1268 ( .A(n1747), .B(n1774), .S(n452), .Z(n1245) );
  MUX2_X1 U1269 ( .A(n1245), .B(n1244), .S(n507), .Z(n1246) );
  MUX2_X1 U1270 ( .A(n1770), .B(n607), .S(n452), .Z(n1247) );
  MUX2_X1 U1271 ( .A(n1805), .B(n603), .S(n452), .Z(n1248) );
  MUX2_X1 U1272 ( .A(n1248), .B(n1247), .S(n507), .Z(n1249) );
  MUX2_X1 U1273 ( .A(n1249), .B(n1246), .S(n1546), .Z(n1250) );
  MUX2_X1 U1274 ( .A(n612), .B(n1753), .S(n452), .Z(n1251) );
  MUX2_X1 U1275 ( .A(n1852), .B(n611), .S(n452), .Z(n1252) );
  MUX2_X1 U1276 ( .A(n1252), .B(n1251), .S(n506), .Z(n1253) );
  MUX2_X1 U1277 ( .A(n1835), .B(n559), .S(n452), .Z(n1254) );
  MUX2_X1 U1278 ( .A(n528), .B(n491), .S(n452), .Z(n1255) );
  MUX2_X1 U1279 ( .A(n526), .B(n1255), .S(n432), .Z(n1256) );
  MUX2_X1 U1280 ( .A(n1256), .B(n1254), .S(n506), .Z(n1257) );
  MUX2_X1 U1281 ( .A(n1257), .B(n1253), .S(n1546), .Z(n1258) );
  MUX2_X1 U1282 ( .A(n1258), .B(n1250), .S(n1566), .Z(n1259) );
  MUX2_X1 U1283 ( .A(n1259), .B(n1243), .S(n1576), .Z(d[36]) );
  MUX2_X1 U1284 ( .A(n1841), .B(n1752), .S(n1548), .Z(n1260) );
  MUX2_X1 U1285 ( .A(n1827), .B(n625), .S(n1546), .Z(n1261) );
  MUX2_X1 U1286 ( .A(n1261), .B(n1260), .S(n507), .Z(n1262) );
  MUX2_X1 U1287 ( .A(n554), .B(n1794), .S(n1546), .Z(n1263) );
  MUX2_X1 U1288 ( .A(n1756), .B(n1772), .S(n1546), .Z(n1264) );
  MUX2_X1 U1289 ( .A(n1264), .B(n1263), .S(n506), .Z(n1265) );
  MUX2_X1 U1290 ( .A(n1265), .B(n1262), .S(n452), .Z(n1266) );
  MUX2_X1 U1291 ( .A(n1767), .B(n1805), .S(n1546), .Z(n1267) );
  MUX2_X1 U1292 ( .A(n1742), .B(n520), .S(n1546), .Z(n1268) );
  MUX2_X1 U1293 ( .A(n1268), .B(n1267), .S(n506), .Z(n1269) );
  MUX2_X1 U1294 ( .A(n1786), .B(n1828), .S(n1547), .Z(n1270) );
  MUX2_X1 U1295 ( .A(n1854), .B(n560), .S(n1547), .Z(n1271) );
  MUX2_X1 U1296 ( .A(n1271), .B(n1270), .S(n508), .Z(n1272) );
  MUX2_X1 U1297 ( .A(n1272), .B(n1269), .S(n453), .Z(n1273) );
  MUX2_X1 U1298 ( .A(n1273), .B(n1266), .S(n1565), .Z(n1274) );
  MUX2_X1 U1299 ( .A(n612), .B(n1758), .S(n1547), .Z(n1275) );
  MUX2_X1 U1301 ( .A(n1276), .B(n1275), .S(n510), .Z(n1277) );
  MUX2_X1 U1302 ( .A(n4870), .B(n552), .S(n1547), .Z(n1278) );
  MUX2_X1 U1303 ( .A(n1842), .B(n1832), .S(n1547), .Z(n1279) );
  MUX2_X1 U1304 ( .A(n1279), .B(n1278), .S(n510), .Z(n1280) );
  MUX2_X1 U1305 ( .A(n1280), .B(n1277), .S(n453), .Z(n1281) );
  MUX2_X1 U1306 ( .A(n1852), .B(n1855), .S(n1547), .Z(n1282) );
  MUX2_X1 U1307 ( .A(n579), .B(n1754), .S(n1547), .Z(n1283) );
  MUX2_X1 U1308 ( .A(n1283), .B(n1282), .S(n510), .Z(n1284) );
  MUX2_X1 U1309 ( .A(n1751), .B(n609), .S(n1547), .Z(n1285) );
  MUX2_X1 U1311 ( .A(n1286), .B(n1285), .S(n510), .Z(n1287) );
  MUX2_X1 U1312 ( .A(n1287), .B(n1284), .S(n453), .Z(n1288) );
  MUX2_X1 U1313 ( .A(n1288), .B(n1281), .S(n1566), .Z(n1289) );
  MUX2_X1 U1314 ( .A(n1289), .B(n1274), .S(n1576), .Z(d[37]) );
  MUX2_X1 U1315 ( .A(n1793), .B(n621), .S(n510), .Z(n1290) );
  MUX2_X1 U1317 ( .A(n1291), .B(n1290), .S(n453), .Z(n1292) );
  MUX2_X1 U1318 ( .A(n1766), .B(n1816), .S(n511), .Z(n1293) );
  MUX2_X1 U1320 ( .A(n1293), .B(n1294), .S(n453), .Z(n1296) );
  MUX2_X1 U1321 ( .A(n1296), .B(n1292), .S(n1547), .Z(n1297) );
  MUX2_X1 U1322 ( .A(n1786), .B(n537), .S(n515), .Z(n1298) );
  MUX2_X1 U1324 ( .A(n1299), .B(n1298), .S(n453), .Z(n1301) );
  MUX2_X1 U1325 ( .A(n622), .B(n593), .S(n511), .Z(n1302) );
  MUX2_X1 U1326 ( .A(n1672), .B(n1302), .S(n453), .Z(n1303) );
  MUX2_X1 U1327 ( .A(n1303), .B(n1301), .S(n1547), .Z(n1304) );
  MUX2_X1 U1328 ( .A(n1304), .B(n1297), .S(n1565), .Z(n1305) );
  MUX2_X1 U1329 ( .A(n579), .B(n578), .S(n511), .Z(n1306) );
  MUX2_X1 U1331 ( .A(n1306), .B(n1307), .S(n453), .Z(n1308) );
  MUX2_X1 U1332 ( .A(n558), .B(n1782), .S(n511), .Z(n1309) );
  MUX2_X1 U1334 ( .A(n1309), .B(n1310), .S(n453), .Z(n1311) );
  MUX2_X1 U1335 ( .A(n1311), .B(n1308), .S(n1547), .Z(n1312) );
  MUX2_X1 U1336 ( .A(n1822), .B(n584), .S(n511), .Z(n1313) );
  MUX2_X1 U1337 ( .A(n629), .B(n612), .S(n511), .Z(n1314) );
  MUX2_X1 U1338 ( .A(n1314), .B(n1313), .S(n453), .Z(n1315) );
  MUX2_X1 U1339 ( .A(n1842), .B(n1799), .S(n511), .Z(n1316) );
  MUX2_X1 U1340 ( .A(n578), .B(n445), .S(n511), .Z(n1317) );
  MUX2_X1 U1341 ( .A(n1317), .B(n1316), .S(n453), .Z(n13180) );
  MUX2_X1 U1342 ( .A(n13180), .B(n1315), .S(n1547), .Z(n1319) );
  MUX2_X1 U1343 ( .A(n1319), .B(n1312), .S(n1566), .Z(n1320) );
  MUX2_X1 U1344 ( .A(n1320), .B(n1305), .S(n1576), .Z(d[38]) );
  MUX2_X1 U1345 ( .A(n595), .B(n1748), .S(n453), .Z(n1321) );
  MUX2_X1 U1347 ( .A(n1321), .B(n1322), .S(n511), .Z(n1323) );
  MUX2_X1 U1348 ( .A(n626), .B(n605), .S(n453), .Z(n1324) );
  MUX2_X1 U1350 ( .A(n1325), .B(n1324), .S(n511), .Z(n1326) );
  MUX2_X1 U1351 ( .A(n1326), .B(n1323), .S(n1547), .Z(n1327) );
  MUX2_X1 U1352 ( .A(n1756), .B(n501), .S(n453), .Z(n1328) );
  MUX2_X1 U1353 ( .A(n1819), .B(n1841), .S(n453), .Z(n1329) );
  MUX2_X1 U1354 ( .A(n1329), .B(n1328), .S(n511), .Z(n1330) );
  MUX2_X1 U1355 ( .A(n570), .B(n1829), .S(n453), .Z(n1331) );
  MUX2_X1 U1356 ( .A(n625), .B(n529), .S(n453), .Z(n1332) );
  MUX2_X1 U1357 ( .A(n1332), .B(n1331), .S(n511), .Z(n13330) );
  MUX2_X1 U1358 ( .A(n13330), .B(n1330), .S(n1547), .Z(n1334) );
  MUX2_X1 U1359 ( .A(n1334), .B(n1327), .S(n1565), .Z(n1335) );
  MUX2_X1 U1360 ( .A(n1769), .B(n1796), .S(n453), .Z(n1336) );
  MUX2_X1 U1362 ( .A(n1337), .B(n1336), .S(n511), .Z(n1338) );
  MUX2_X1 U1363 ( .A(n527), .B(n1807), .S(n454), .Z(n1339) );
  MUX2_X1 U1364 ( .A(n552), .B(n618), .S(n454), .Z(n1340) );
  MUX2_X1 U1365 ( .A(n1340), .B(n1339), .S(n511), .Z(n1341) );
  MUX2_X1 U1366 ( .A(n1341), .B(n1338), .S(n1547), .Z(n1342) );
  MUX2_X1 U1367 ( .A(n1845), .B(n1826), .S(n454), .Z(n1343) );
  MUX2_X1 U1368 ( .A(n1757), .B(n1343), .S(n511), .Z(n1344) );
  MUX2_X1 U1369 ( .A(n1827), .B(n1745), .S(n457), .Z(n1345) );
  MUX2_X1 U1370 ( .A(n598), .B(n540), .S(n454), .Z(n1346) );
  MUX2_X1 U1371 ( .A(n1346), .B(n1345), .S(n511), .Z(n1347) );
  MUX2_X1 U1372 ( .A(n1347), .B(n1344), .S(n1547), .Z(n1348) );
  MUX2_X1 U1373 ( .A(n1348), .B(n1342), .S(n1565), .Z(n1349) );
  MUX2_X1 U1374 ( .A(n1349), .B(n1335), .S(n1576), .Z(d[39]) );
  MUX2_X1 U1375 ( .A(n611), .B(n1776), .S(n454), .Z(n1350) );
  MUX2_X1 U1376 ( .A(n1754), .B(n1745), .S(n454), .Z(n1351) );
  MUX2_X1 U1377 ( .A(n1351), .B(n1350), .S(n511), .Z(n13520) );
  MUX2_X1 U1379 ( .A(n13520), .B(n1353), .S(n1547), .Z(n1355) );
  MUX2_X1 U1380 ( .A(n547), .B(n1746), .S(n454), .Z(n1356) );
  MUX2_X1 U1381 ( .A(n1813), .B(n1674), .S(n454), .Z(n1357) );
  MUX2_X1 U1382 ( .A(n1357), .B(n1356), .S(n511), .Z(n1358) );
  MUX2_X1 U1383 ( .A(n1834), .B(n620), .S(n454), .Z(n1359) );
  MUX2_X1 U1384 ( .A(n1814), .B(n550), .S(n454), .Z(n1360) );
  MUX2_X1 U1385 ( .A(n1360), .B(n1359), .S(n512), .Z(n1361) );
  MUX2_X1 U1386 ( .A(n1361), .B(n1358), .S(n1547), .Z(n1362) );
  MUX2_X1 U1387 ( .A(n1362), .B(n1355), .S(n1565), .Z(n1363) );
  MUX2_X1 U1388 ( .A(n1805), .B(n1808), .S(n454), .Z(n1364) );
  MUX2_X1 U1390 ( .A(n1365), .B(n1364), .S(n512), .Z(n1367) );
  MUX2_X1 U1391 ( .A(n1746), .B(n605), .S(n454), .Z(n1368) );
  MUX2_X1 U1393 ( .A(n593), .B(n1369), .S(n454), .Z(n1370) );
  MUX2_X1 U1394 ( .A(n1370), .B(n1368), .S(n512), .Z(n1371) );
  MUX2_X1 U1395 ( .A(n1371), .B(n1367), .S(addr[5]), .Z(n1372) );
  MUX2_X1 U1396 ( .A(n569), .B(n561), .S(n454), .Z(n1373) );
  MUX2_X1 U1397 ( .A(n1810), .B(n1751), .S(n454), .Z(n1374) );
  MUX2_X1 U1398 ( .A(n1374), .B(n1373), .S(n512), .Z(n1375) );
  MUX2_X1 U1399 ( .A(n562), .B(n1776), .S(n454), .Z(n1376) );
  MUX2_X1 U1400 ( .A(n523), .B(n620), .S(n454), .Z(n1377) );
  MUX2_X1 U1401 ( .A(n1377), .B(n1376), .S(n512), .Z(n1378) );
  MUX2_X1 U1402 ( .A(n1378), .B(n1375), .S(addr[5]), .Z(n1379) );
  MUX2_X1 U1403 ( .A(n1379), .B(n1372), .S(n1565), .Z(n1380) );
  MUX2_X1 U1404 ( .A(n1380), .B(n1363), .S(n1576), .Z(d[3]) );
  MUX2_X1 U1405 ( .A(n618), .B(n1813), .S(n455), .Z(n1381) );
  MUX2_X1 U1406 ( .A(n543), .B(n1802), .S(n455), .Z(n1382) );
  MUX2_X1 U1407 ( .A(n1382), .B(n1381), .S(n512), .Z(n1383) );
  MUX2_X1 U1408 ( .A(n578), .B(n616), .S(n455), .Z(n1384) );
  MUX2_X1 U1409 ( .A(n528), .B(n520), .S(n455), .Z(n1385) );
  MUX2_X1 U1410 ( .A(n1385), .B(n1384), .S(n512), .Z(n1386) );
  MUX2_X1 U1411 ( .A(n1386), .B(n1383), .S(n1543), .Z(n1387) );
  MUX2_X1 U1412 ( .A(n1771), .B(n1829), .S(n455), .Z(n1388) );
  MUX2_X1 U1413 ( .A(n543), .B(n1756), .S(n455), .Z(n1389) );
  MUX2_X1 U1414 ( .A(n1389), .B(n1388), .S(n512), .Z(n1390) );
  MUX2_X1 U1415 ( .A(n548), .B(n1774), .S(n455), .Z(n1391) );
  MUX2_X1 U1416 ( .A(n586), .B(n599), .S(n455), .Z(n1392) );
  MUX2_X1 U1417 ( .A(n1392), .B(n1391), .S(n512), .Z(n1393) );
  MUX2_X1 U1418 ( .A(n1393), .B(n1390), .S(addr[5]), .Z(n1394) );
  MUX2_X1 U1419 ( .A(n1394), .B(n1387), .S(n1565), .Z(n1395) );
  MUX2_X1 U1420 ( .A(n526), .B(n1765), .S(n455), .Z(n1396) );
  MUX2_X1 U1421 ( .A(n611), .B(n581), .S(n455), .Z(n1397) );
  MUX2_X1 U1422 ( .A(n1397), .B(n1396), .S(n512), .Z(n1398) );
  MUX2_X1 U1423 ( .A(n564), .B(n596), .S(n455), .Z(n1399) );
  MUX2_X1 U1424 ( .A(n608), .B(n1813), .S(n455), .Z(n1400) );
  MUX2_X1 U1425 ( .A(n1400), .B(n1399), .S(n512), .Z(n1401) );
  MUX2_X1 U1426 ( .A(n1401), .B(n1398), .S(addr[5]), .Z(n1402) );
  MUX2_X1 U1427 ( .A(n1797), .B(n1801), .S(n512), .Z(n1403) );
  MUX2_X1 U1428 ( .A(n1850), .B(n1403), .S(n428), .Z(n1404) );
  MUX2_X1 U1429 ( .A(n526), .B(n601), .S(n455), .Z(n1405) );
  MUX2_X1 U1431 ( .A(n1406), .B(n1405), .S(n512), .Z(n1407) );
  MUX2_X1 U1432 ( .A(n1407), .B(n1404), .S(addr[5]), .Z(n1408) );
  MUX2_X1 U1433 ( .A(n1408), .B(n1402), .S(n1565), .Z(n1409) );
  MUX2_X1 U1434 ( .A(n1409), .B(n1395), .S(n1576), .Z(d[40]) );
  MUX2_X1 U1435 ( .A(n536), .B(n621), .S(n512), .Z(n1410) );
  MUX2_X1 U1437 ( .A(n1411), .B(n1410), .S(n455), .Z(n1412) );
  MUX2_X1 U1438 ( .A(n444), .B(n1854), .S(n512), .Z(n1413) );
  MUX2_X1 U1439 ( .A(n1830), .B(n564), .S(n512), .Z(n1414) );
  MUX2_X1 U1440 ( .A(n1414), .B(n1413), .S(n455), .Z(n1415) );
  MUX2_X1 U1441 ( .A(n1415), .B(n1412), .S(n1548), .Z(n1416) );
  MUX2_X1 U1442 ( .A(addr[0]), .B(n590), .S(n512), .Z(n1417) );
  MUX2_X1 U1443 ( .A(n1832), .B(n1761), .S(n512), .Z(n1418) );
  MUX2_X1 U1444 ( .A(n1418), .B(n1417), .S(n455), .Z(n1419) );
  MUX2_X1 U1445 ( .A(n517), .B(n1850), .S(n513), .Z(n1420) );
  MUX2_X1 U1446 ( .A(n1752), .B(n621), .S(n513), .Z(n1421) );
  MUX2_X1 U1447 ( .A(n1421), .B(n1420), .S(n455), .Z(n1422) );
  MUX2_X1 U1448 ( .A(n1422), .B(n1419), .S(addr[5]), .Z(n1423) );
  MUX2_X1 U1449 ( .A(n1423), .B(n1416), .S(n1565), .Z(n1424) );
  MUX2_X1 U1450 ( .A(n1761), .B(n601), .S(n513), .Z(n1425) );
  MUX2_X1 U1451 ( .A(n595), .B(addr[0]), .S(n513), .Z(n1426) );
  MUX2_X1 U1452 ( .A(n1426), .B(n1425), .S(n455), .Z(n1427) );
  MUX2_X1 U1453 ( .A(n535), .B(n575), .S(n513), .Z(n1428) );
  MUX2_X1 U1455 ( .A(n1428), .B(n1429), .S(n456), .Z(n1430) );
  MUX2_X1 U1456 ( .A(n1430), .B(n1427), .S(addr[5]), .Z(n1431) );
  MUX2_X1 U1457 ( .A(n760), .B(n611), .S(n513), .Z(n1432) );
  MUX2_X1 U1458 ( .A(n1830), .B(n1766), .S(n513), .Z(n1433) );
  MUX2_X1 U1459 ( .A(n1433), .B(n1432), .S(n456), .Z(n1434) );
  MUX2_X1 U1460 ( .A(n531), .B(n1815), .S(n513), .Z(n1435) );
  MUX2_X1 U1461 ( .A(n1793), .B(n605), .S(n513), .Z(n1436) );
  MUX2_X1 U1462 ( .A(n1436), .B(n1435), .S(n456), .Z(n1437) );
  MUX2_X1 U1463 ( .A(n1437), .B(n1434), .S(addr[5]), .Z(n1438) );
  MUX2_X1 U1464 ( .A(n1438), .B(n1431), .S(n1565), .Z(n1439) );
  MUX2_X1 U1465 ( .A(n1439), .B(n1424), .S(n1576), .Z(d[41]) );
  MUX2_X1 U1466 ( .A(n1809), .B(n1794), .S(n513), .Z(n1440) );
  MUX2_X1 U1467 ( .A(addr[0]), .B(n585), .S(n513), .Z(n1441) );
  MUX2_X1 U1468 ( .A(n1441), .B(n1440), .S(n456), .Z(n1442) );
  MUX2_X1 U1469 ( .A(n4870), .B(n554), .S(n513), .Z(n1443) );
  MUX2_X1 U1470 ( .A(n584), .B(n1833), .S(n513), .Z(n1444) );
  MUX2_X1 U1471 ( .A(n1444), .B(n1443), .S(n456), .Z(n1445) );
  MUX2_X1 U1472 ( .A(n1445), .B(n1442), .S(n1545), .Z(n1446) );
  MUX2_X1 U1473 ( .A(n443), .B(n530), .S(n513), .Z(n1447) );
  MUX2_X1 U1475 ( .A(n1448), .B(n1447), .S(n456), .Z(n1449) );
  MUX2_X1 U1476 ( .A(n1844), .B(n1764), .S(n513), .Z(n1450) );
  MUX2_X1 U1477 ( .A(n530), .B(n618), .S(n513), .Z(n1451) );
  MUX2_X1 U1478 ( .A(n1451), .B(n1450), .S(n456), .Z(n1452) );
  MUX2_X1 U1479 ( .A(n1452), .B(n1449), .S(n1549), .Z(n1453) );
  MUX2_X1 U1480 ( .A(n1453), .B(n1446), .S(n1565), .Z(n1454) );
  MUX2_X1 U1481 ( .A(n1773), .B(n612), .S(n513), .Z(n1455) );
  MUX2_X1 U1482 ( .A(n1797), .B(n445), .S(n513), .Z(n1456) );
  MUX2_X1 U1483 ( .A(n1456), .B(n1455), .S(n456), .Z(n1457) );
  MUX2_X1 U1484 ( .A(n526), .B(n612), .S(n514), .Z(n1458) );
  MUX2_X1 U1485 ( .A(n1458), .B(n633), .S(n456), .Z(n1459) );
  MUX2_X1 U1486 ( .A(n1459), .B(n1457), .S(addr[5]), .Z(n1460) );
  MUX2_X1 U1487 ( .A(n1750), .B(n540), .S(n514), .Z(n1461) );
  MUX2_X1 U1488 ( .A(n1832), .B(n593), .S(n514), .Z(n1462) );
  MUX2_X1 U1489 ( .A(n1462), .B(n1461), .S(n456), .Z(n1463) );
  MUX2_X1 U1490 ( .A(n523), .B(n1852), .S(n514), .Z(n1464) );
  MUX2_X1 U1491 ( .A(n545), .B(n1847), .S(n514), .Z(n1465) );
  MUX2_X1 U1492 ( .A(n1465), .B(n1464), .S(n456), .Z(n1466) );
  MUX2_X1 U1493 ( .A(n1466), .B(n1463), .S(addr[5]), .Z(n1467) );
  MUX2_X1 U1494 ( .A(n1467), .B(n1460), .S(n1565), .Z(n1468) );
  MUX2_X1 U1495 ( .A(n1468), .B(n1454), .S(n1576), .Z(d[42]) );
  MUX2_X1 U1496 ( .A(n4870), .B(n501), .S(n514), .Z(n1469) );
  MUX2_X1 U1497 ( .A(n1469), .B(n1673), .S(n456), .Z(n1470) );
  MUX2_X1 U1498 ( .A(n579), .B(n1764), .S(n514), .Z(n1471) );
  MUX2_X1 U1499 ( .A(n533), .B(n1786), .S(n514), .Z(n1472) );
  MUX2_X1 U1500 ( .A(n1472), .B(n1471), .S(n456), .Z(n1473) );
  MUX2_X1 U1501 ( .A(n1473), .B(n1470), .S(n1550), .Z(n1474) );
  MUX2_X1 U1502 ( .A(n444), .B(n567), .S(n514), .Z(n1475) );
  MUX2_X1 U1503 ( .A(n535), .B(n1829), .S(n514), .Z(n1476) );
  MUX2_X1 U1504 ( .A(n1476), .B(n1475), .S(n456), .Z(n1477) );
  MUX2_X1 U1505 ( .A(n1755), .B(n612), .S(n514), .Z(n1478) );
  MUX2_X1 U1506 ( .A(n1773), .B(n493), .S(n514), .Z(n1479) );
  MUX2_X1 U1507 ( .A(n1479), .B(n1478), .S(n456), .Z(n1480) );
  MUX2_X1 U1508 ( .A(n1480), .B(n1477), .S(n1551), .Z(n1481) );
  MUX2_X1 U1509 ( .A(n1481), .B(n1474), .S(n1565), .Z(n1482) );
  MUX2_X1 U1510 ( .A(n1798), .B(n564), .S(n514), .Z(n1483) );
  MUX2_X1 U1511 ( .A(n1787), .B(addr[2]), .S(n514), .Z(n1484) );
  MUX2_X1 U1512 ( .A(n1484), .B(n1483), .S(n456), .Z(n1485) );
  MUX2_X1 U1513 ( .A(n1843), .B(n502), .S(n514), .Z(n1486) );
  MUX2_X1 U1514 ( .A(n1673), .B(n1486), .S(n456), .Z(n1487) );
  MUX2_X1 U1515 ( .A(n1487), .B(n1485), .S(addr[5]), .Z(n1488) );
  MUX2_X1 U1516 ( .A(n1761), .B(n1764), .S(n514), .Z(n1489) );
  MUX2_X1 U1517 ( .A(n563), .B(n1802), .S(n514), .Z(n1490) );
  MUX2_X1 U1518 ( .A(n1490), .B(n1489), .S(n456), .Z(n1491) );
  MUX2_X1 U1519 ( .A(n553), .B(n577), .S(n514), .Z(n1492) );
  MUX2_X1 U1520 ( .A(n1811), .B(n605), .S(n515), .Z(n1493) );
  MUX2_X1 U1521 ( .A(n1493), .B(n1492), .S(n457), .Z(n1494) );
  MUX2_X1 U1522 ( .A(n1494), .B(n1491), .S(addr[5]), .Z(n1495) );
  MUX2_X1 U1523 ( .A(n1495), .B(n1488), .S(n1565), .Z(n1496) );
  MUX2_X1 U1524 ( .A(n1496), .B(n1482), .S(n1576), .Z(d[43]) );
  XOR2_X1 U1525 ( .A(n615), .B(n506), .Z(n1070) );
  MUX2_X1 U1526 ( .A(n528), .B(n502), .S(n432), .Z(n1497) );
  MUX2_X1 U1537 ( .A(addr[0]), .B(n1498), .S(n1548), .Z(n1502) );
  MUX2_X1 U1538 ( .A(n627), .B(n1792), .S(n515), .Z(n1503) );
  MUX2_X1 U1539 ( .A(addr[0]), .B(n525), .S(n515), .Z(n734) );
  MUX2_X1 U1540 ( .A(n445), .B(n1794), .S(n515), .Z(n1504) );
  MUX2_X1 U1541 ( .A(n1782), .B(n1816), .S(n457), .Z(n765) );
  MUX2_X1 U1542 ( .A(n500), .B(n1843), .S(n432), .Z(n1505) );
  MUX2_X1 U1543 ( .A(n526), .B(n4870), .S(n432), .Z(n1506) );
  MUX2_X1 U1544 ( .A(n1840), .B(n572), .S(n457), .Z(n855) );
  MUX2_X1 U1545 ( .A(n1820), .B(n628), .S(n457), .Z(n884) );
  MUX2_X1 U1546 ( .A(addr[2]), .B(n502), .S(n433), .Z(n1507) );
  MUX2_X1 U1547 ( .A(n604), .B(n1807), .S(n457), .Z(n1508) );
  MUX2_X1 U1548 ( .A(n4870), .B(n1800), .S(n432), .Z(n1509) );
  MUX2_X1 U1549 ( .A(n526), .B(n517), .S(n432), .Z(n1510) );
  MUX2_X1 U1550 ( .A(n560), .B(n1809), .S(n457), .Z(n1027) );
  MUX2_X1 U1551 ( .A(addr[2]), .B(n1760), .S(n515), .Z(n1511) );
  MUX2_X1 U1552 ( .A(n628), .B(n1837), .S(n457), .Z(n1084) );
  MUX2_X1 U1553 ( .A(n1750), .B(n1829), .S(n432), .Z(n1512) );
  MUX2_X1 U1554 ( .A(n444), .B(n593), .S(n515), .Z(n1513) );
  MUX2_X1 U1556 ( .A(n1513), .B(n1514), .S(n1545), .Z(n1116) );
  MUX2_X1 U1557 ( .A(n1843), .B(n502), .S(n432), .Z(n1515) );
  MUX2_X1 U1558 ( .A(n1505), .B(n1765), .S(n457), .Z(n1160) );
  MUX2_X1 U1559 ( .A(addr[2]), .B(n1829), .S(n432), .Z(n1516) );
  MUX2_X1 U1560 ( .A(n1809), .B(n1758), .S(n457), .Z(n1517) );
  MUX2_X1 U1561 ( .A(n501), .B(n517), .S(n432), .Z(n1518) );
  MUX2_X1 U1562 ( .A(n1763), .B(n1804), .S(n457), .Z(n1354) );
  MUX2_X1 U1563 ( .A(n520), .B(n528), .S(n450), .Z(n1366) );
  MUX2_X1 U1564 ( .A(n629), .B(n593), .S(n515), .Z(n1519) );
  DFF_X1 c1_reg_17_ ( .D(n409), .CK(clk), .Q(c1[17]) );
  NAND2_X1 U3 ( .A1(n1664), .A2(n408), .ZN(n409) );
  INV_X1 U4 ( .A(n1688), .ZN(n408) );
  INV_X1 U5 ( .A(n518), .ZN(n1756) );
  INV_X1 U6 ( .A(n558), .ZN(n1773) );
  INV_X1 U7 ( .A(n48), .ZN(n1611) );
  INV_X1 U8 ( .A(n538), .ZN(n1755) );
  INV_X1 U9 ( .A(n27), .ZN(n1607) );
  INV_X1 U10 ( .A(n520), .ZN(n1829) );
  INV_X1 U11 ( .A(n9), .ZN(n1858) );
  INV_X1 U12 ( .A(n6), .ZN(n1861) );
  NAND2_X1 U13 ( .A1(n9), .A2(n10), .ZN(n8) );
  INV_X1 U14 ( .A(n2), .ZN(n1857) );
  INV_X1 U17 ( .A(n627), .ZN(n1802) );
  NAND2_X1 U18 ( .A1(n520), .A2(n543), .ZN(n542) );
  NAND2_X1 U20 ( .A1(n450), .A2(n1701), .ZN(n1694) );
  NAND2_X1 U22 ( .A1(n543), .A2(n1782), .ZN(n558) );
  INV_X1 U28 ( .A(n529), .ZN(n1821) );
  NAND2_X1 U30 ( .A1(n519), .A2(n520), .ZN(n518) );
  NAND2_X1 U37 ( .A1(n519), .A2(n1782), .ZN(n538) );
  NAND2_X1 U39 ( .A1(n7), .A2(n2), .ZN(n27) );
  INV_X1 U44 ( .A(n525), .ZN(n1810) );
  INV_X1 U46 ( .A(n628), .ZN(n1830) );
  INV_X1 U47 ( .A(n531), .ZN(n1837) );
  INV_X1 U49 ( .A(n583), .ZN(n1786) );
  AOI21_X1 U53 ( .B1(n450), .B2(n587), .A(n609), .ZN(n1337) );
  NAND2_X1 U55 ( .A1(n6), .A2(n4), .ZN(n48) );
  INV_X1 U56 ( .A(n524), .ZN(n1820) );
  INV_X1 U58 ( .A(n565), .ZN(n1788) );
  NAND2_X1 U106 ( .A1(n6), .A2(n10), .ZN(n15) );
  NAND2_X1 U130 ( .A1(n2), .A2(n4), .ZN(n261) );
  INV_X1 U147 ( .A(n537), .ZN(n1793) );
  INV_X1 U168 ( .A(n58), .ZN(n1643) );
  INV_X1 U170 ( .A(n1708), .ZN(n1856) );
  NAND2_X1 U191 ( .A1(n450), .A2(n1745), .ZN(n1230) );
  NAND2_X1 U192 ( .A1(n450), .A2(n529), .ZN(n742) );
  INV_X1 U196 ( .A(n609), .ZN(n1745) );
  INV_X1 U201 ( .A(n563), .ZN(n1764) );
  INV_X1 U203 ( .A(n590), .ZN(n1761) );
  INV_X1 U205 ( .A(n532), .ZN(n1791) );
  INV_X1 U206 ( .A(n589), .ZN(n1797) );
  INV_X1 U208 ( .A(n552), .ZN(n1754) );
  INV_X1 U213 ( .A(n571), .ZN(n1776) );
  INV_X1 U223 ( .A(n588), .ZN(n1805) );
  INV_X1 U248 ( .A(n619), .ZN(n1826) );
  INV_X1 U252 ( .A(n587), .ZN(n1743) );
  INV_X1 U259 ( .A(n548), .ZN(n1769) );
  INV_X1 U261 ( .A(n559), .ZN(n1765) );
  INV_X1 U262 ( .A(n578), .ZN(n1832) );
  INV_X1 U268 ( .A(n527), .ZN(n1811) );
  INV_X1 U300 ( .A(n557), .ZN(n1789) );
  INV_X1 U309 ( .A(n560), .ZN(n1808) );
  INV_X1 U313 ( .A(n585), .ZN(n1742) );
  INV_X1 U318 ( .A(n10), .ZN(n1646) );
  INV_X1 U329 ( .A(n550), .ZN(n1790) );
  INV_X1 U344 ( .A(n530), .ZN(n1771) );
  INV_X1 U348 ( .A(n620), .ZN(n1841) );
  INV_X1 U352 ( .A(n564), .ZN(n1775) );
  INV_X1 U355 ( .A(n547), .ZN(n1833) );
  INV_X1 U359 ( .A(n626), .ZN(n1844) );
  INV_X1 U381 ( .A(n4), .ZN(n1610) );
  INV_X1 U403 ( .A(n605), .ZN(n1778) );
  INV_X1 U408 ( .A(n603), .ZN(n1759) );
  INV_X1 U409 ( .A(n31), .ZN(n1625) );
  INV_X1 U410 ( .A(n553), .ZN(n1674) );
  INV_X1 U411 ( .A(n541), .ZN(n1767) );
  INV_X1 U412 ( .A(n204), .ZN(n1650) );
  INV_X1 U413 ( .A(n606), .ZN(n1779) );
  NOR2_X1 U414 ( .A1(n1782), .A2(n1837), .ZN(n410) );
  INV_X1 U415 ( .A(n625), .ZN(n1758) );
  AND3_X1 U416 ( .A1(n1858), .A2(n4), .A3(n248), .ZN(n247) );
  INV_X1 U417 ( .A(n522), .ZN(n1770) );
  INV_X1 U418 ( .A(n584), .ZN(n1741) );
  INV_X1 U419 ( .A(n598), .ZN(n1850) );
  INV_X1 U437 ( .A(n572), .ZN(n1796) );
  INV_X1 U440 ( .A(n566), .ZN(n1795) );
  INV_X1 U441 ( .A(n19), .ZN(n1614) );
  INV_X1 U442 ( .A(n575), .ZN(n1763) );
  INV_X1 U443 ( .A(n596), .ZN(n1824) );
  INV_X1 U444 ( .A(n26), .ZN(n1622) );
  INV_X1 U445 ( .A(n43), .ZN(n1634) );
  INV_X1 U446 ( .A(n750), .ZN(n1669) );
  INV_X1 U447 ( .A(n545), .ZN(n1766) );
  INV_X1 U448 ( .A(n21), .ZN(n1617) );
  INV_X1 U449 ( .A(n556), .ZN(n1835) );
  INV_X1 U450 ( .A(n622), .ZN(n1827) );
  INV_X1 U451 ( .A(n576), .ZN(n1839) );
  INV_X1 U452 ( .A(n49), .ZN(n1638) );
  INV_X1 U453 ( .A(n582), .ZN(n1838) );
  INV_X1 U454 ( .A(n51), .ZN(n1640) );
  NAND2_X1 U455 ( .A1(n1836), .A2(n1295), .ZN(n1294) );
  INV_X1 U456 ( .A(n542), .ZN(n1836) );
  NAND2_X1 U457 ( .A1(n1633), .A2(n248), .ZN(n354) );
  INV_X1 U458 ( .A(n570), .ZN(n1846) );
  INV_X1 U459 ( .A(n595), .ZN(n1804) );
  INV_X1 U460 ( .A(n591), .ZN(n1777) );
  INV_X1 U461 ( .A(n22), .ZN(n1618) );
  INV_X1 U462 ( .A(n32), .ZN(n1626) );
  INV_X1 U463 ( .A(n56), .ZN(n1641) );
  INV_X1 U464 ( .A(n610), .ZN(n1784) );
  INV_X1 U465 ( .A(n611), .ZN(n1831) );
  INV_X1 U466 ( .A(n3), .ZN(n1612) );
  INV_X1 U467 ( .A(n613), .ZN(n1845) );
  INV_X1 U468 ( .A(n221), .ZN(n1645) );
  INV_X1 U469 ( .A(n20), .ZN(n1616) );
  INV_X1 U470 ( .A(n47), .ZN(n1637) );
  INV_X1 U471 ( .A(n50), .ZN(n1639) );
  INV_X1 U472 ( .A(n24), .ZN(n1620) );
  INV_X1 U473 ( .A(n34), .ZN(n1628) );
  INV_X1 U474 ( .A(n607), .ZN(n1840) );
  AND2_X1 U475 ( .A1(n1300), .A2(n519), .ZN(n1307) );
  INV_X1 U476 ( .A(n1517), .ZN(n1757) );
  INV_X1 U477 ( .A(n18), .ZN(n1613) );
  INV_X1 U478 ( .A(n39), .ZN(n1630) );
  INV_X1 U479 ( .A(n1680), .ZN(n1664) );
  NAND2_X1 U480 ( .A1(addr[2]), .A2(addr[3]), .ZN(n520) );
  INV_X1 U481 ( .A(n533), .ZN(n1782) );
  NAND2_X1 U482 ( .A1(n432), .A2(n4640), .ZN(n2) );
  INV_X1 U483 ( .A(n476), .ZN(n452) );
  INV_X1 U484 ( .A(n478), .ZN(n457) );
  INV_X1 U485 ( .A(n475), .ZN(n450) );
  INV_X1 U486 ( .A(n475), .ZN(n449) );
  INV_X1 U487 ( .A(n475), .ZN(n463) );
  NOR2_X1 U488 ( .A1(addr[3]), .A2(n485), .ZN(n1701) );
  NAND2_X1 U489 ( .A1(n435), .A2(n526), .ZN(n525) );
  NAND2_X1 U490 ( .A1(n533), .A2(n525), .ZN(n532) );
  INV_X1 U491 ( .A(n5), .ZN(n1859) );
  NAND2_X1 U492 ( .A1(n435), .A2(n449), .ZN(n6) );
  NAND2_X1 U493 ( .A1(n432), .A2(n520), .ZN(n531) );
  INV_X1 U494 ( .A(n517), .ZN(n1750) );
  NAND2_X1 U495 ( .A1(n433), .A2(n517), .ZN(n519) );
  NAND2_X1 U496 ( .A1(n485), .A2(n466), .ZN(n1708) );
  INV_X1 U497 ( .A(n528), .ZN(n1843) );
  INV_X1 U498 ( .A(n526), .ZN(n1800) );
  NAND2_X1 U499 ( .A1(n433), .A2(n528), .ZN(n543) );
  NAND2_X1 U500 ( .A1(n1543), .A2(n1), .ZN(n4) );
  NAND2_X1 U501 ( .A1(n434), .A2(n1782), .ZN(n522) );
  NAND2_X1 U502 ( .A1(addr[0]), .A2(n1829), .ZN(n529) );
  NAND2_X1 U503 ( .A1(n1544), .A2(n504), .ZN(n1680) );
  INV_X1 U504 ( .A(n1), .ZN(n1860) );
  NAND2_X1 U505 ( .A1(n517), .A2(n522), .ZN(n523) );
  XNOR2_X1 U506 ( .A(n5), .B(n1545), .ZN(n411) );
  NAND2_X1 U507 ( .A1(n521), .A2(n520), .ZN(n548) );
  NAND2_X1 U508 ( .A1(n1544), .A2(n5), .ZN(n10) );
  NAND2_X1 U509 ( .A1(n528), .A2(n525), .ZN(n527) );
  OAI21_X1 U510 ( .B1(n1700), .B2(n1701), .A(n1589), .ZN(n1676) );
  NOR2_X1 U511 ( .A1(addr[3]), .A2(n1859), .ZN(n1700) );
  NAND2_X1 U512 ( .A1(n543), .A2(n517), .ZN(n625) );
  INV_X1 U513 ( .A(n551), .ZN(n1792) );
  NOR2_X1 U514 ( .A1(addr[3]), .A2(n1856), .ZN(n1693) );
  NOR2_X1 U515 ( .A1(addr[3]), .A2(n434), .ZN(n1726) );
  NAND2_X1 U516 ( .A1(addr[0]), .A2(n1800), .ZN(n537) );
  NAND2_X1 U517 ( .A1(n517), .A2(n531), .ZN(n541) );
  NAND2_X1 U518 ( .A1(n517), .A2(n525), .ZN(n545) );
  NAND2_X1 U519 ( .A1(n531), .A2(n526), .ZN(n560) );
  NOR2_X1 U520 ( .A1(n469), .A2(n485), .ZN(n1685) );
  INV_X1 U521 ( .A(n539), .ZN(n1794) );
  NAND2_X1 U522 ( .A1(n6), .A2(n1543), .ZN(n19) );
  NAND2_X1 U523 ( .A1(addr[0]), .A2(addr[3]), .ZN(n524) );
  NAND2_X1 U524 ( .A1(n1544), .A2(n1857), .ZN(n130) );
  NAND2_X1 U525 ( .A1(n522), .A2(n528), .ZN(n530) );
  NAND2_X1 U526 ( .A1(n1544), .A2(n1858), .ZN(n7) );
  NAND2_X1 U527 ( .A1(n434), .A2(n1750), .ZN(n587) );
  NAND2_X1 U528 ( .A1(n528), .A2(n519), .ZN(n552) );
  NAND2_X1 U529 ( .A1(n1543), .A2(n1860), .ZN(n21) );
  NAND2_X1 U530 ( .A1(n1701), .A2(n1702), .ZN(n1690) );
  NAND2_X1 U531 ( .A1(n519), .A2(n526), .ZN(n760) );
  INV_X1 U532 ( .A(n536), .ZN(n1809) );
  NAND2_X1 U533 ( .A1(n1544), .A2(n2), .ZN(n58) );
  INV_X1 U534 ( .A(n569), .ZN(n1834) );
  NAND2_X1 U535 ( .A1(n526), .A2(n543), .ZN(n776) );
  NAND2_X1 U536 ( .A1(n505), .A2(n558), .ZN(n1295) );
  NAND2_X1 U537 ( .A1(n1579), .A2(n55), .ZN(n248) );
  NAND2_X1 U538 ( .A1(n531), .A2(n528), .ZN(n582) );
  NAND2_X1 U539 ( .A1(n4), .A2(n5), .ZN(n3) );
  OR2_X1 U540 ( .A1(n1858), .A2(n1552), .ZN(n13) );
  NAND2_X1 U541 ( .A1(n505), .A2(n1821), .ZN(n750) );
  INV_X1 U542 ( .A(n1684), .ZN(n1589) );
  NAND2_X1 U543 ( .A1(n1544), .A2(n1861), .ZN(n46) );
  AOI21_X1 U544 ( .B1(n449), .B2(n616), .A(n1786), .ZN(n1204) );
  NAND2_X1 U545 ( .A1(n58), .A2(n5), .ZN(n57) );
  INV_X1 U546 ( .A(n561), .ZN(n1774) );
  NAND2_X1 U547 ( .A1(n505), .A2(n563), .ZN(n1300) );
  OAI21_X1 U548 ( .B1(n1687), .B2(n1688), .A(n1689), .ZN(n1678) );
  NAND3_X1 U549 ( .A1(n1586), .A2(n1690), .A3(n504), .ZN(n1689) );
  AOI21_X1 U550 ( .B1(n1543), .B2(n565), .A(n1794), .ZN(n1276) );
  NAND2_X1 U551 ( .A1(n471), .A2(n1543), .ZN(n204) );
  AOI21_X1 U552 ( .B1(n1578), .B2(n53), .A(n17), .ZN(n252) );
  INV_X1 U553 ( .A(n54), .ZN(n1615) );
  INV_X1 U555 ( .A(n629), .ZN(n1854) );
  NAND2_X1 U558 ( .A1(n5), .A2(n19), .ZN(n105) );
  AOI21_X1 U559 ( .B1(n505), .B2(n571), .A(n1816), .ZN(n1024) );
  AOI21_X1 U560 ( .B1(n505), .B2(n527), .A(n1765), .ZN(n869) );
  AOI21_X1 U561 ( .B1(n449), .B2(n561), .A(n1743), .ZN(n1166) );
  NAND2_X1 U562 ( .A1(n1859), .A2(n1543), .ZN(n43) );
  INV_X1 U565 ( .A(n579), .ZN(n1812) );
  INV_X1 U568 ( .A(n535), .ZN(n1823) );
  INV_X1 U570 ( .A(n616), .ZN(n1783) );
  NAND2_X1 U579 ( .A1(n1), .A2(n19), .ZN(n54) );
  INV_X1 U585 ( .A(n593), .ZN(n1813) );
  INV_X1 U591 ( .A(n417), .ZN(n1598) );
  NOR2_X1 U592 ( .A1(n504), .A2(n1051), .ZN(n1055) );
  NOR2_X1 U593 ( .A1(addr[3]), .A2(n1859), .ZN(n198) );
  NOR2_X1 U598 ( .A1(n1564), .A2(n1810), .ZN(n710) );
  NOR2_X1 U603 ( .A1(n1577), .A2(n522), .ZN(n993) );
  NOR2_X1 U604 ( .A1(n1578), .A2(n28), .ZN(n351) );
  NAND2_X1 U608 ( .A1(n505), .A2(n1823), .ZN(n1110) );
  NAND2_X1 U611 ( .A1(n1843), .A2(n434), .ZN(n607) );
  INV_X1 U615 ( .A(n1511), .ZN(n1672) );
  INV_X1 U618 ( .A(n422), .ZN(n1659) );
  INV_X1 U627 ( .A(n1519), .ZN(n1673) );
  INV_X1 U635 ( .A(n1502), .ZN(n1663) );
  INV_X1 U636 ( .A(n414), .ZN(n1652) );
  INV_X1 U646 ( .A(n418), .ZN(n1655) );
  INV_X1 U649 ( .A(n419), .ZN(n1656) );
  INV_X1 U671 ( .A(n415), .ZN(n1653) );
  INV_X1 U677 ( .A(n44), .ZN(n1635) );
  INV_X1 U687 ( .A(n416), .ZN(n1654) );
  INV_X1 U702 ( .A(n1510), .ZN(n1752) );
  OAI21_X1 U705 ( .B1(n1849), .B2(n467), .A(n524), .ZN(n1325) );
  INV_X1 U707 ( .A(n567), .ZN(n1807) );
  INV_X1 U724 ( .A(n581), .ZN(n1849) );
  AOI21_X1 U726 ( .B1(addr[3]), .B2(n311), .A(n1599), .ZN(n310) );
  INV_X1 U728 ( .A(n55), .ZN(n1600) );
  AOI21_X1 U731 ( .B1(addr[3]), .B2(n23), .A(n1661), .ZN(n298) );
  NAND2_X1 U747 ( .A1(n402), .A2(n403), .ZN(n401) );
  INV_X1 U748 ( .A(n8), .ZN(n1648) );
  INV_X1 U750 ( .A(n41), .ZN(n1632) );
  INV_X1 U754 ( .A(n35), .ZN(n1595) );
  INV_X1 U756 ( .A(n38), .ZN(n1597) );
  INV_X1 U757 ( .A(n1706), .ZN(n1590) );
  OAI21_X1 U765 ( .B1(n1543), .B2(n1687), .A(n1564), .ZN(n1706) );
  INV_X1 U773 ( .A(n601), .ZN(n1798) );
  INV_X1 U775 ( .A(n586), .ZN(n1762) );
  INV_X1 U779 ( .A(n555), .ZN(n1855) );
  NOR2_X1 U790 ( .A1(n469), .A2(n569), .ZN(n743) );
  INV_X1 U809 ( .A(n554), .ZN(n1772) );
  INV_X1 U811 ( .A(n29), .ZN(n1594) );
  INV_X1 U822 ( .A(n612), .ZN(n1803) );
  INV_X1 U831 ( .A(n604), .ZN(n1853) );
  INV_X1 U838 ( .A(n42), .ZN(n1633) );
  OAI21_X1 U840 ( .B1(n1108), .B2(n1109), .A(n1116), .ZN(n1115) );
  NAND2_X1 U851 ( .A1(n535), .A2(n1295), .ZN(n1448) );
  INV_X1 U858 ( .A(n11), .ZN(n1591) );
  AOI21_X1 U869 ( .B1(n505), .B2(n13), .A(n1643), .ZN(n379) );
  AOI21_X1 U883 ( .B1(n347), .B2(n1577), .A(n341), .ZN(n346) );
  NAND2_X1 U887 ( .A1(n521), .A2(n526), .ZN(n1369) );
  NOR2_X1 U898 ( .A1(n504), .A2(n936), .ZN(n940) );
  NOR2_X1 U911 ( .A1(n504), .A2(n965), .ZN(n969) );
  NOR2_X1 U925 ( .A1(n1543), .A2(n534), .ZN(n694) );
  NOR2_X1 U927 ( .A1(n504), .A2(n1810), .ZN(n692) );
  INV_X1 U947 ( .A(n817), .ZN(n1781) );
  INV_X1 U956 ( .A(n540), .ZN(n1847) );
  INV_X1 U984 ( .A(n25), .ZN(n1621) );
  INV_X1 U986 ( .A(n17), .ZN(n1609) );
  INV_X1 U1011 ( .A(n407), .ZN(n1603) );
  INV_X1 U1012 ( .A(n13), .ZN(n1608) );
  INV_X1 U1015 ( .A(n57), .ZN(n1644) );
  INV_X1 U1043 ( .A(n59), .ZN(n1642) );
  NOR2_X1 U1045 ( .A1(n1564), .A2(n1790), .ZN(n794) );
  INV_X1 U1074 ( .A(n608), .ZN(n1785) );
  OAI21_X1 U1080 ( .B1(n470), .B2(n579), .A(n593), .ZN(n932) );
  AOI21_X1 U1102 ( .B1(n1543), .B2(n536), .A(n1752), .ZN(n1286) );
  AOI21_X1 U1104 ( .B1(n449), .B2(n627), .A(n585), .ZN(n1406) );
  NOR2_X1 U1112 ( .A1(n485), .A2(n1650), .ZN(n168) );
  NOR2_X1 U1129 ( .A1(n1564), .A2(n533), .ZN(n638) );
  NOR2_X1 U1131 ( .A1(n1564), .A2(n517), .ZN(n844) );
  AND2_X1 U1134 ( .A1(n578), .A2(n474), .ZN(n1086) );
  AOI21_X1 U1152 ( .B1(n223), .B2(addr[3]), .A(n220), .ZN(n222) );
  NOR2_X1 U1156 ( .A1(n1188), .A2(n1186), .ZN(n1200) );
  NAND2_X1 U1158 ( .A1(n434), .A2(n465), .ZN(n736) );
  INV_X1 U1162 ( .A(n519), .ZN(n1753) );
  NOR2_X1 U1179 ( .A1(n1860), .A2(n1643), .ZN(n358) );
  INV_X1 U1185 ( .A(n16), .ZN(n1593) );
  NOR2_X1 U1190 ( .A1(n600), .A2(n821), .ZN(n825) );
  NOR2_X1 U1207 ( .A1(n1577), .A2(n1744), .ZN(n997) );
  INV_X1 U1210 ( .A(n406), .ZN(n1602) );
  INV_X1 U1212 ( .A(n23), .ZN(n1619) );
  INV_X1 U1220 ( .A(n7), .ZN(n1606) );
  INV_X1 U1225 ( .A(n15), .ZN(n1647) );
  NAND2_X1 U1228 ( .A1(n2), .A2(n10), .ZN(n328) );
  NOR2_X1 U1252 ( .A1(n1543), .A2(n1859), .ZN(n342) );
  INV_X1 U1253 ( .A(n562), .ZN(n1848) );
  NOR2_X1 U1300 ( .A1(n1564), .A2(n1802), .ZN(n635) );
  NOR2_X1 U1310 ( .A1(n504), .A2(n908), .ZN(n912) );
  NAND2_X1 U1316 ( .A1(n1853), .A2(n449), .ZN(n910) );
  NOR2_X1 U1319 ( .A1(n504), .A2(n1794), .ZN(n1094) );
  INV_X1 U1323 ( .A(n546), .ZN(n1585) );
  NOR2_X1 U1330 ( .A1(n537), .A2(n4680), .ZN(n1229) );
  AOI21_X1 U1333 ( .B1(n504), .B2(n529), .A(n626), .ZN(n1310) );
  AND2_X1 U1346 ( .A1(n585), .A2(n474), .ZN(n1322) );
  NAND2_X1 U1349 ( .A1(n505), .A2(n588), .ZN(n1411) );
  OAI21_X1 U1361 ( .B1(n470), .B2(n589), .A(n525), .ZN(n1171) );
  NAND2_X1 U1378 ( .A1(n1366), .A2(n525), .ZN(n1365) );
  NAND2_X1 U1389 ( .A1(n734), .A2(n465), .ZN(n733) );
  NOR2_X1 U1392 ( .A1(n504), .A2(n731), .ZN(n732) );
  INV_X1 U1430 ( .A(n33), .ZN(n1627) );
  INV_X1 U1436 ( .A(n594), .ZN(n1760) );
  OR2_X1 U1454 ( .A1(n1685), .A2(n1565), .ZN(n1683) );
  INV_X1 U1474 ( .A(n36), .ZN(n1596) );
  INV_X1 U1527 ( .A(n311), .ZN(n1605) );
  INV_X1 U1528 ( .A(n573), .ZN(n1787) );
  INV_X1 U1529 ( .A(n592), .ZN(n1744) );
  INV_X1 U1530 ( .A(n614), .ZN(n1825) );
  INV_X1 U1531 ( .A(n544), .ZN(n1852) );
  INV_X1 U1532 ( .A(n602), .ZN(n1815) );
  INV_X1 U1533 ( .A(n837), .ZN(n1842) );
  INV_X1 U1534 ( .A(n424), .ZN(n1661) );
  INV_X1 U1535 ( .A(n599), .ZN(n1814) );
  INV_X1 U1536 ( .A(n40), .ZN(n1631) );
  INV_X1 U1555 ( .A(n617), .ZN(n1746) );
  INV_X1 U1565 ( .A(n615), .ZN(n1780) );
  INV_X1 U1566 ( .A(n632), .ZN(n1667) );
  INV_X1 U1567 ( .A(n618), .ZN(n1747) );
  INV_X1 U1568 ( .A(n621), .ZN(n1748) );
  INV_X1 U1569 ( .A(n130), .ZN(n1649) );
  NAND2_X1 U1570 ( .A1(n1635), .A2(n317), .ZN(n316) );
  OAI21_X1 U1571 ( .B1(n430), .B2(n1861), .A(addr[3]), .ZN(n317) );
  INV_X1 U1572 ( .A(n1498), .ZN(n1668) );
  INV_X1 U1573 ( .A(n521), .ZN(n1768) );
  INV_X1 U1574 ( .A(n549), .ZN(n1822) );
  INV_X1 U1575 ( .A(n1505), .ZN(n1817) );
  INV_X1 U1576 ( .A(n37), .ZN(n1629) );
  AND2_X1 U1577 ( .A1(n1300), .A2(n837), .ZN(n1299) );
  INV_X1 U1578 ( .A(n425), .ZN(n1662) );
  INV_X1 U1579 ( .A(n421), .ZN(n1658) );
  INV_X1 U1580 ( .A(n423), .ZN(n1660) );
  INV_X1 U1581 ( .A(n412), .ZN(n1604) );
  INV_X1 U1582 ( .A(n28), .ZN(n1623) );
  INV_X1 U1583 ( .A(n1503), .ZN(n1670) );
  INV_X1 U1584 ( .A(n1516), .ZN(n1828) );
  INV_X1 U1585 ( .A(n420), .ZN(n1657) );
  INV_X1 U1586 ( .A(n1512), .ZN(n1749) );
  INV_X1 U1587 ( .A(n1508), .ZN(n1806) );
  INV_X1 U1588 ( .A(n46), .ZN(n1636) );
  INV_X1 U1589 ( .A(n30), .ZN(n1624) );
  INV_X1 U1590 ( .A(n479), .ZN(n460) );
  INV_X1 U1591 ( .A(n477), .ZN(n454) );
  INV_X1 U1592 ( .A(n479), .ZN(n461) );
  INV_X1 U1593 ( .A(n474), .ZN(n462) );
  INV_X1 U1594 ( .A(n476), .ZN(n451) );
  INV_X1 U1595 ( .A(n477), .ZN(n455) );
  INV_X1 U1596 ( .A(n478), .ZN(n456) );
  INV_X1 U1597 ( .A(n479), .ZN(n459) );
  INV_X1 U1598 ( .A(n477), .ZN(n453) );
  INV_X1 U1599 ( .A(n476), .ZN(n458) );
  NOR2_X1 U1600 ( .A1(n1543), .A2(n1564), .ZN(n1699) );
  OAI21_X1 U1601 ( .B1(n1565), .B2(n485), .A(n1684), .ZN(n1729) );
  NAND2_X1 U1602 ( .A1(addr[3]), .A2(n504), .ZN(n1682) );
  NAND2_X1 U1603 ( .A1(n1579), .A2(n1564), .ZN(n1688) );
  INV_X1 U1604 ( .A(n12), .ZN(n1592) );
  NOR2_X1 U1605 ( .A1(n1680), .A2(n1704), .ZN(n1697) );
  INV_X1 U1606 ( .A(n1704), .ZN(n1586) );
  NAND2_X1 U1607 ( .A1(addr[3]), .A2(n1592), .ZN(n189) );
  INV_X1 U1608 ( .A(n52), .ZN(n1599) );
  AND2_X1 U1609 ( .A1(n1697), .A2(n435), .ZN(n1728) );
  NAND2_X1 U1610 ( .A1(n1544), .A2(n1666), .ZN(n1187) );
  INV_X1 U1611 ( .A(n624), .ZN(n1666) );
  NAND2_X1 U1612 ( .A1(n482), .A2(n494), .ZN(n517) );
  NAND2_X1 U1613 ( .A1(n497), .A2(n486), .ZN(n526) );
  NAND2_X1 U1614 ( .A1(addr[3]), .A2(n486), .ZN(n528) );
  INV_X1 U1615 ( .A(n1536), .ZN(n504) );
  INV_X1 U1616 ( .A(n1560), .ZN(n1543) );
  INV_X1 U1617 ( .A(n1536), .ZN(n506) );
  INV_X1 U1618 ( .A(n1560), .ZN(n1545) );
  INV_X1 U1619 ( .A(n500), .ZN(n489) );
  INV_X1 U1620 ( .A(n437), .ZN(n435) );
  INV_X1 U1621 ( .A(n1536), .ZN(n505) );
  INV_X1 U1622 ( .A(n1537), .ZN(n5090) );
  INV_X1 U1623 ( .A(n1560), .ZN(n1548) );
  INV_X1 U1624 ( .A(n1538), .ZN(n513) );
  INV_X1 U1625 ( .A(n1537), .ZN(n514) );
  INV_X1 U1626 ( .A(n1538), .ZN(n515) );
  INV_X1 U1627 ( .A(n1538), .ZN(n1521) );
  INV_X1 U1628 ( .A(n1539), .ZN(n1522) );
  INV_X1 U1629 ( .A(n1539), .ZN(n1523) );
  INV_X1 U1630 ( .A(n1539), .ZN(n1524) );
  INV_X1 U1631 ( .A(n1537), .ZN(n510) );
  INV_X1 U1632 ( .A(n1538), .ZN(n1500) );
  INV_X1 U1633 ( .A(n1537), .ZN(n512) );
  INV_X1 U1634 ( .A(n1537), .ZN(n511) );
  INV_X1 U1635 ( .A(n1539), .ZN(n1501) );
  INV_X1 U1636 ( .A(n1539), .ZN(n1520) );
  INV_X1 U1637 ( .A(n1537), .ZN(n508) );
  INV_X1 U1638 ( .A(n1538), .ZN(n516) );
  INV_X1 U1639 ( .A(n1560), .ZN(n1551) );
  INV_X1 U1640 ( .A(n1538), .ZN(n1499) );
  INV_X1 U1641 ( .A(n1536), .ZN(n507) );
  INV_X1 U1642 ( .A(n442), .ZN(n433) );
  INV_X1 U1643 ( .A(n1561), .ZN(n1550) );
  INV_X1 U1644 ( .A(n1561), .ZN(n1549) );
  INV_X1 U1645 ( .A(n443), .ZN(n434) );
  INV_X1 U1646 ( .A(n1583), .ZN(n1579) );
  INV_X1 U1647 ( .A(n1583), .ZN(n1578) );
  INV_X1 U1648 ( .A(n497), .ZN(n493) );
  INV_X1 U1649 ( .A(n442), .ZN(n432) );
  NAND2_X1 U1650 ( .A1(n471), .A2(n438), .ZN(n5) );
  INV_X1 U1651 ( .A(n1559), .ZN(n1544) );
  NAND2_X1 U1652 ( .A1(n533), .A2(n436), .ZN(n616) );
  NAND2_X1 U1653 ( .A1(n441), .A2(n449), .ZN(n1) );
  AOI221_X1 U1654 ( .B1(n408), .B2(n1680), .C1(n1699), .C2(n1720), .A(n1721), 
        .ZN(n1719) );
  NOR3_X1 U1655 ( .A1(n1582), .A2(n1564), .A3(n1859), .ZN(n1721) );
  OAI221_X1 U1656 ( .B1(n1722), .B2(n1708), .C1(n1723), .C2(n1531), .A(n1724), 
        .ZN(n1720) );
  NAND2_X1 U1657 ( .A1(n1544), .A2(n1569), .ZN(n1684) );
  INV_X1 U1658 ( .A(n1559), .ZN(n1552) );
  NAND2_X1 U1659 ( .A1(n441), .A2(n526), .ZN(n536) );
  NAND2_X1 U1660 ( .A1(addr[0]), .A2(n494), .ZN(n593) );
  NAND2_X1 U1661 ( .A1(n483), .A2(n439), .ZN(n555) );
  AOI221_X1 U1662 ( .B1(n1713), .B2(n1699), .C1(n1532), .C2(n1589), .A(n1714), 
        .ZN(n1712) );
  AOI21_X1 U1663 ( .B1(n1715), .B2(n1684), .A(n435), .ZN(n1714) );
  OAI21_X1 U1664 ( .B1(n1680), .B2(n1701), .A(n1564), .ZN(n1715) );
  NAND2_X1 U1665 ( .A1(n1829), .A2(n438), .ZN(n535) );
  NAND2_X1 U1666 ( .A1(n520), .A2(n437), .ZN(n569) );
  OAI221_X1 U1667 ( .B1(n1543), .B2(n1730), .C1(n1664), .C2(n1581), .A(n1731), 
        .ZN(N1333) );
  AOI21_X1 U1668 ( .B1(n1735), .B2(n1525), .A(n1736), .ZN(n1730) );
  NOR3_X1 U1669 ( .A1(n1732), .A2(n1586), .A3(n1733), .ZN(n1731) );
  NOR3_X1 U1670 ( .A1(n4680), .A2(n1726), .A3(n1528), .ZN(n1736) );
  OAI221_X1 U1671 ( .B1(n1578), .B2(n1675), .C1(n1534), .C2(n1676), .A(n1677), 
        .ZN(N509) );
  AOI22_X1 U1672 ( .A1(n1678), .A2(n1553), .B1(n1579), .B2(n1679), .ZN(n1677)
         );
  AOI22_X1 U1673 ( .A1(n1543), .A2(n1691), .B1(n1692), .B2(n1569), .ZN(n1675)
         );
  OAI221_X1 U1674 ( .B1(n1680), .B2(n1681), .C1(n1682), .C2(n1683), .A(n1684), 
        .ZN(n1679) );
  OAI221_X1 U1675 ( .B1(n1590), .B2(n1582), .C1(n506), .C2(n1684), .A(n1696), 
        .ZN(N487) );
  AOI221_X1 U1676 ( .B1(n1697), .B2(n1690), .C1(n1698), .C2(n1699), .A(n1588), 
        .ZN(n1696) );
  AND2_X1 U1677 ( .A1(n1694), .A2(n505), .ZN(n1698) );
  INV_X1 U1678 ( .A(n1676), .ZN(n1588) );
  NAND2_X1 U1679 ( .A1(n442), .A2(n1800), .ZN(n539) );
  NAND2_X1 U1680 ( .A1(n493), .A2(n439), .ZN(n581) );
  OAI22_X1 U1681 ( .A1(n505), .A2(n1693), .B1(n1532), .B2(n1694), .ZN(n1692)
         );
  NAND2_X1 U1682 ( .A1(n450), .A2(n1555), .ZN(n38) );
  NAND2_X1 U1683 ( .A1(n441), .A2(n528), .ZN(n540) );
  NAND2_X1 U1684 ( .A1(n498), .A2(n439), .ZN(n551) );
  NAND2_X1 U1685 ( .A1(n1859), .A2(n1554), .ZN(n36) );
  AOI22_X1 U1686 ( .A1(n1725), .A2(n4640), .B1(n1726), .B2(n449), .ZN(n1723)
         );
  OAI21_X1 U1687 ( .B1(n1579), .B2(n494), .A(n440), .ZN(n1725) );
  NAND2_X1 U1688 ( .A1(n520), .A2(n1526), .ZN(n574) );
  NAND2_X1 U1689 ( .A1(n442), .A2(n517), .ZN(n897) );
  NAND2_X1 U1690 ( .A1(n433), .A2(n1556), .ZN(n311) );
  OAI21_X1 U1691 ( .B1(n1533), .B2(n1837), .A(n535), .ZN(n534) );
  OAI21_X1 U1692 ( .B1(n505), .B2(n1685), .A(n1587), .ZN(n1691) );
  INV_X1 U1693 ( .A(n1695), .ZN(n1587) );
  AOI21_X1 U1694 ( .B1(n1690), .B2(n504), .A(n1570), .ZN(n1695) );
  NAND2_X1 U1695 ( .A1(n1782), .A2(n438), .ZN(n817) );
  NAND2_X1 U1696 ( .A1(n2), .A2(n1554), .ZN(n29) );
  AOI21_X1 U1697 ( .B1(n1694), .B2(n1734), .A(n505), .ZN(n1732) );
  NAND3_X1 U1698 ( .A1(n473), .A2(n496), .A3(n432), .ZN(n1734) );
  AOI21_X1 U1699 ( .B1(n1762), .B2(n1569), .A(n1533), .ZN(n600) );
  OAI21_X1 U1700 ( .B1(n628), .B2(n1570), .A(n577), .ZN(n717) );
  NAND2_X1 U1701 ( .A1(n434), .A2(n486), .ZN(n544) );
  NAND2_X1 U1702 ( .A1(n5), .A2(n486), .ZN(n45) );
  NAND2_X1 U1703 ( .A1(n1693), .A2(n1526), .ZN(n1687) );
  NAND2_X1 U1704 ( .A1(n1843), .A2(n436), .ZN(n837) );
  NAND2_X1 U1705 ( .A1(n472), .A2(n437), .ZN(n1702) );
  OAI21_X1 U1706 ( .B1(n1686), .B2(n1856), .A(n496), .ZN(n1681) );
  NOR2_X1 U1707 ( .A1(n435), .A2(n486), .ZN(n1686) );
  OR2_X1 U1708 ( .A1(n1782), .A2(n443), .ZN(n521) );
  NAND4_X1 U1709 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .ZN(N1352)
         );
  OAI211_X1 U1710 ( .C1(n1544), .C2(n1713), .A(n1586), .B(n449), .ZN(n1716) );
  NAND4_X1 U1711 ( .A1(n1859), .A2(n1729), .A3(n1525), .A4(n1580), .ZN(n1717)
         );
  OAI211_X1 U1712 ( .C1(n1727), .C2(n1728), .A(n484), .B(addr[3]), .ZN(n1718)
         );
  NAND2_X1 U1713 ( .A1(n497), .A2(n204), .ZN(n203) );
  AOI21_X1 U1714 ( .B1(addr[3]), .B2(n36), .A(n18), .ZN(n205) );
  AOI21_X1 U1715 ( .B1(n493), .B2(n11), .A(n29), .ZN(n306) );
  NAND2_X1 U1716 ( .A1(n1860), .A2(n1555), .ZN(n55) );
  NAND2_X1 U1717 ( .A1(n1557), .A2(n1861), .ZN(n11) );
  AOI21_X1 U1718 ( .B1(n1709), .B2(n1710), .A(n1577), .ZN(N1975) );
  NAND4_X1 U1719 ( .A1(n1699), .A2(n449), .A3(n1711), .A4(n436), .ZN(n1710) );
  OR2_X1 U1720 ( .A1(n1712), .A2(n463), .ZN(n1709) );
  OAI22_X1 U1721 ( .A1(addr[3]), .A2(n1528), .B1(n505), .B2(n1701), .ZN(n1711)
         );
  OAI211_X1 U1722 ( .C1(n1590), .C2(n1582), .A(n1703), .B(n1704), .ZN(N468) );
  OAI211_X1 U1723 ( .C1(n1705), .C2(n489), .A(n1581), .B(n1664), .ZN(n1703) );
  NOR2_X1 U1724 ( .A1(n486), .A2(n1702), .ZN(n1705) );
  NAND2_X1 U1725 ( .A1(n1858), .A2(n1556), .ZN(n406) );
  NAND2_X1 U1726 ( .A1(n1), .A2(n1555), .ZN(n407) );
  NAND2_X1 U1727 ( .A1(n1750), .A2(n440), .ZN(n592) );
  NAND2_X1 U1728 ( .A1(n505), .A2(n21), .ZN(n426) );
  NAND2_X1 U1729 ( .A1(n486), .A2(n440), .ZN(n604) );
  AND2_X1 U1730 ( .A1(n6), .A2(n1556), .ZN(n427) );
  INV_X1 U1731 ( .A(n1507), .ZN(n1818) );
  INV_X1 U1732 ( .A(n1504), .ZN(n1671) );
  INV_X1 U1733 ( .A(n1509), .ZN(n1799) );
  INV_X1 U1734 ( .A(n1518), .ZN(n1751) );
  NAND2_X1 U1735 ( .A1(n1823), .A2(n1527), .ZN(n1514) );
  OAI21_X1 U1736 ( .B1(n497), .B2(n1601), .A(n130), .ZN(n129) );
  INV_X1 U1737 ( .A(n62), .ZN(n1601) );
  OAI21_X1 U1738 ( .B1(n1534), .B2(n1794), .A(n1783), .ZN(n967) );
  OAI21_X1 U1739 ( .B1(n1792), .B2(n1529), .A(n593), .ZN(n873) );
  OAI21_X1 U1740 ( .B1(n13), .B2(n495), .A(n36), .ZN(n211) );
  OAI21_X1 U1741 ( .B1(n1788), .B2(n1529), .A(n1774), .ZN(n1061) );
  OAI21_X1 U1742 ( .B1(n1571), .B2(n1821), .A(n1771), .ZN(n807) );
  OAI21_X1 U1743 ( .B1(n1571), .B2(n1802), .A(n817), .ZN(n816) );
  OAI21_X1 U1744 ( .B1(n1582), .B2(n1643), .A(n130), .ZN(n267) );
  OAI21_X1 U1745 ( .B1(n1582), .B2(n48), .A(n53), .ZN(n259) );
  OAI21_X1 U1746 ( .B1(n1778), .B2(n1581), .A(n539), .ZN(n994) );
  OAI21_X1 U1747 ( .B1(n1646), .B2(n495), .A(n12), .ZN(n193) );
  NAND2_X1 U1748 ( .A1(n1558), .A2(n1857), .ZN(n16) );
  NAND2_X1 U1749 ( .A1(n1582), .A2(n547), .ZN(n546) );
  NOR2_X1 U1750 ( .A1(addr[3]), .A2(n1557), .ZN(n188) );
  AND2_X1 U1751 ( .A1(n201), .A2(n1572), .ZN(n200) );
  NOR2_X1 U1752 ( .A1(n1707), .A2(n1688), .ZN(N464) );
  AOI22_X1 U1753 ( .A1(n1687), .A2(n1553), .B1(n1544), .B2(n1682), .ZN(n1707)
         );
  NAND2_X1 U1754 ( .A1(n1834), .A2(n1526), .ZN(n1498) );
  XNOR2_X1 U1755 ( .A(n1535), .B(n450), .ZN(n428) );
  NOR2_X1 U1756 ( .A1(n568), .A2(n664), .ZN(n665) );
  NOR2_X1 U1757 ( .A1(n1821), .A2(n1581), .ZN(n1133) );
  NOR2_X1 U1758 ( .A1(n791), .A2(n792), .ZN(n796) );
  NOR2_X1 U1759 ( .A1(n548), .A2(n1570), .ZN(n597) );
  XNOR2_X1 U1760 ( .A(n498), .B(n484), .ZN(n429) );
  INV_X1 U1761 ( .A(n1497), .ZN(n1816) );
  OAI21_X1 U1762 ( .B1(n1849), .B2(n1530), .A(n551), .ZN(n1429) );
  AND2_X1 U1763 ( .A1(n855), .A2(n1535), .ZN(n854) );
  OAI22_X1 U1764 ( .A1(n1532), .A2(n580), .B1(n1834), .B2(n467), .ZN(n740) );
  NOR2_X1 U1765 ( .A1(n1809), .A2(n449), .ZN(n580) );
  NOR2_X1 U1766 ( .A1(n432), .A2(n1564), .ZN(n714) );
  AOI21_X1 U1767 ( .B1(n1564), .B2(n759), .A(n450), .ZN(n758) );
  OAI22_X1 U1768 ( .A1(n525), .A2(n1528), .B1(n1668), .B2(n1557), .ZN(n759) );
  OAI21_X1 U1769 ( .B1(n1571), .B2(n565), .A(n837), .ZN(n836) );
  NOR2_X1 U1770 ( .A1(n1793), .A2(n1530), .ZN(n689) );
  INV_X1 U1771 ( .A(n574), .ZN(n1665) );
  NOR2_X1 U1772 ( .A1(n536), .A2(n1531), .ZN(n1112) );
  OAI22_X1 U1773 ( .A1(n431), .A2(n466), .B1(n1578), .B2(n435), .ZN(n1139) );
  NAND2_X1 U1774 ( .A1(n551), .A2(n1580), .ZN(n1137) );
  NOR2_X1 U1775 ( .A1(n1861), .A2(n486), .ZN(n146) );
  OAI21_X1 U1776 ( .B1(n1533), .B2(n566), .A(n565), .ZN(n675) );
  AND2_X1 U1777 ( .A1(n765), .A2(n1532), .ZN(n764) );
  AND2_X1 U1778 ( .A1(n884), .A2(n1533), .ZN(n883) );
  AND2_X1 U1779 ( .A1(n1027), .A2(n1536), .ZN(n1026) );
  NOR2_X1 U1780 ( .A1(n449), .A2(n1669), .ZN(n1192) );
  NAND2_X1 U1781 ( .A1(n1792), .A2(n1527), .ZN(n1190) );
  AND2_X1 U1782 ( .A1(n1354), .A2(n1535), .ZN(n1353) );
  NOR2_X1 U1783 ( .A1(n1858), .A2(n1561), .ZN(n430) );
  AND2_X1 U1784 ( .A1(n433), .A2(n1580), .ZN(n431) );
  NAND2_X1 U1785 ( .A1(n1792), .A2(n1580), .ZN(n1143) );
  AND2_X1 U1786 ( .A1(n523), .A2(n1572), .ZN(n660) );
  AND2_X1 U1787 ( .A1(n1825), .A2(n1535), .ZN(n1291) );
  AND2_X1 U1788 ( .A1(n1084), .A2(n1535), .ZN(n1083) );
  AND2_X1 U1789 ( .A1(n1160), .A2(n1536), .ZN(n1159) );
  INV_X1 U1790 ( .A(n1506), .ZN(n1801) );
  INV_X1 U1791 ( .A(n413), .ZN(n1651) );
  INV_X1 U1792 ( .A(n1515), .ZN(n1819) );
  NAND2_X1 U1793 ( .A1(n12), .A2(n486), .ZN(n166) );
  INV_X1 U1794 ( .A(n45), .ZN(n1851) );
  INV_X1 U1795 ( .A(n1573), .ZN(n1564) );
  INV_X1 U1796 ( .A(n1560), .ZN(n1546) );
  INV_X1 U1797 ( .A(n1561), .ZN(n1547) );
  INV_X1 U1798 ( .A(n1573), .ZN(n1567) );
  INV_X1 U1799 ( .A(n1573), .ZN(n1566) );
  INV_X1 U1800 ( .A(n499), .ZN(n492) );
  INV_X1 U1801 ( .A(n500), .ZN(n491) );
  INV_X1 U1802 ( .A(n500), .ZN(n490) );
  INV_X1 U1803 ( .A(n1574), .ZN(n1568) );
  INV_X1 U1804 ( .A(n1573), .ZN(n1565) );
  NOR3_X1 U1805 ( .A1(n1684), .A2(n1529), .A3(n1581), .ZN(n1727) );
  NAND2_X1 U1806 ( .A1(n472), .A2(n1553), .ZN(n12) );
  OAI221_X1 U1807 ( .B1(n504), .B2(n1738), .C1(n1544), .C2(n1531), .A(n1739), 
        .ZN(N1318) );
  NOR2_X1 U1808 ( .A1(n1589), .A2(n1586), .ZN(n1739) );
  AOI221_X1 U1809 ( .B1(n449), .B2(n485), .C1(addr[3]), .C2(n1740), .A(n1578), 
        .ZN(n1738) );
  NAND2_X1 U1810 ( .A1(n1859), .A2(n486), .ZN(n1740) );
  NAND2_X1 U1811 ( .A1(n1565), .A2(n1581), .ZN(n1704) );
  NAND3_X1 U1812 ( .A1(n450), .A2(n1530), .A3(addr[3]), .ZN(n1724) );
  AOI21_X1 U1813 ( .B1(n496), .B2(n1580), .A(n435), .ZN(n1722) );
  AOI21_X1 U1814 ( .B1(n1859), .B2(n1525), .A(n1684), .ZN(n1733) );
  OAI21_X1 U1815 ( .B1(addr[3]), .B2(n1708), .A(n1737), .ZN(n1735) );
  NAND3_X1 U1816 ( .A1(addr[3]), .A2(n486), .A3(n1859), .ZN(n1737) );
  NAND2_X1 U1817 ( .A1(n450), .A2(n1527), .ZN(n624) );
  NAND2_X1 U1818 ( .A1(n493), .A2(n1554), .ZN(n14) );
  NOR2_X1 U1819 ( .A1(n1564), .A2(n486), .ZN(n823) );
  NAND2_X1 U1820 ( .A1(n441), .A2(n1682), .ZN(n1713) );
  NAND2_X1 U1821 ( .A1(n1558), .A2(n437), .ZN(n52) );
  NAND3_X1 U1822 ( .A1(n1572), .A2(n495), .A3(n38), .ZN(n207) );
  AND4_X1 U1823 ( .A1(n1583), .A2(n1682), .A3(n1699), .A4(n1859), .ZN(N1952)
         );
  BUF_X1 U1824 ( .A(n1540), .Z(n1538) );
  BUF_X1 U1825 ( .A(n1540), .Z(n1537) );
  BUF_X1 U1826 ( .A(n1542), .Z(n1539) );
  BUF_X1 U1827 ( .A(n1563), .Z(n1560) );
  BUF_X1 U1828 ( .A(n1541), .Z(n1536) );
  BUF_X1 U1829 ( .A(n1563), .Z(n1561) );
  BUF_X1 U1830 ( .A(n447), .Z(n442) );
  BUF_X1 U1831 ( .A(n495), .Z(n500) );
  BUF_X1 U1832 ( .A(n503), .Z(n499) );
  BUF_X1 U1833 ( .A(n1563), .Z(n1559) );
  BUF_X1 U1834 ( .A(n447), .Z(n438) );
  BUF_X1 U1835 ( .A(n447), .Z(n439) );
  BUF_X1 U1836 ( .A(n447), .Z(n437) );
  BUF_X1 U1837 ( .A(n447), .Z(n443) );
  BUF_X1 U1838 ( .A(n494), .Z(n497) );
  BUF_X1 U1839 ( .A(n447), .Z(n436) );
  BUF_X1 U1840 ( .A(n447), .Z(n440) );
  BUF_X1 U1841 ( .A(n447), .Z(n441) );
  BUF_X1 U1842 ( .A(n496), .Z(n501) );
  BUF_X1 U1843 ( .A(n488), .Z(n486) );
  BUF_X1 U1844 ( .A(n503), .Z(n498) );
  BUF_X1 U1845 ( .A(n503), .Z(n494) );
  BUF_X1 U1846 ( .A(n488), .Z(n4870) );
  BUF_X1 U1847 ( .A(n1584), .Z(n1583) );
  BUF_X1 U1848 ( .A(n1584), .Z(n1580) );
  AND3_X1 U1849 ( .A1(n1565), .A2(n1528), .A3(n520), .ZN(n712) );
  BUF_X1 U1850 ( .A(n1575), .Z(n1573) );
  BUF_X1 U1851 ( .A(n447), .Z(n444) );
  BUF_X1 U1852 ( .A(n447), .Z(n445) );
  BUF_X1 U1853 ( .A(n1542), .Z(n1525) );
  BUF_X1 U1854 ( .A(n503), .Z(n495) );
  BUF_X1 U1855 ( .A(n1542), .Z(n1532) );
  BUF_X1 U1856 ( .A(n1542), .Z(n1533) );
  BUF_X1 U1857 ( .A(n1562), .Z(n1558) );
  BUF_X1 U1858 ( .A(n1542), .Z(n1534) );
  BUF_X1 U1859 ( .A(n1554), .Z(n1557) );
  BUF_X1 U1860 ( .A(n503), .Z(n496) );
  BUF_X1 U1861 ( .A(n1575), .Z(n1569) );
  BUF_X1 U1862 ( .A(n1562), .Z(n1553) );
  BUF_X1 U1863 ( .A(n1542), .Z(n1527) );
  BUF_X1 U1864 ( .A(n1542), .Z(n1526) );
  BUF_X1 U1865 ( .A(n1562), .Z(n1554) );
  BUF_X1 U1866 ( .A(n1562), .Z(n1556) );
  BUF_X1 U1867 ( .A(n1562), .Z(n1555) );
  BUF_X1 U1868 ( .A(n1530), .Z(n1528) );
  BUF_X1 U1869 ( .A(n1584), .Z(n1581) );
  BUF_X1 U1870 ( .A(n1541), .Z(n1535) );
  BUF_X1 U1871 ( .A(n1531), .Z(n1529) );
  BUF_X1 U1872 ( .A(n1535), .Z(n1530) );
  BUF_X1 U1873 ( .A(n1542), .Z(n1531) );
  BUF_X1 U1874 ( .A(n1575), .Z(n1570) );
  BUF_X1 U1875 ( .A(n1575), .Z(n1574) );
  BUF_X1 U1876 ( .A(n1584), .Z(n1582) );
  BUF_X1 U1877 ( .A(n1575), .Z(n1572) );
  BUF_X1 U1878 ( .A(n1575), .Z(n1571) );
  BUF_X1 U1879 ( .A(n496), .Z(n502) );
  BUF_X1 U1880 ( .A(n1559), .Z(n1562) );
  BUF_X1 U1881 ( .A(n447), .Z(n446) );
  INV_X1 U1882 ( .A(addr[2]), .ZN(n488) );
  INV_X1 U1883 ( .A(addr[3]), .ZN(n503) );
  INV_X1 U1884 ( .A(addr[7]), .ZN(n1584) );
  INV_X1 U1885 ( .A(addr[0]), .ZN(n447) );
  BUF_X1 U1886 ( .A(addr[1]), .Z(n448) );
  BUF_X1 U1887 ( .A(n481), .Z(n4640) );
  BUF_X1 U1888 ( .A(n470), .Z(n465) );
  BUF_X1 U1889 ( .A(n465), .Z(n466) );
  BUF_X1 U1890 ( .A(n470), .Z(n467) );
  BUF_X1 U1891 ( .A(n469), .Z(n4680) );
  BUF_X1 U1892 ( .A(n480), .Z(n469) );
  BUF_X1 U1893 ( .A(n480), .Z(n470) );
  BUF_X1 U1894 ( .A(n481), .Z(n471) );
  BUF_X1 U1895 ( .A(n4640), .Z(n472) );
  BUF_X1 U1896 ( .A(n481), .Z(n473) );
  BUF_X1 U1897 ( .A(n478), .Z(n474) );
  BUF_X1 U1898 ( .A(n481), .Z(n475) );
  BUF_X1 U1899 ( .A(n472), .Z(n476) );
  BUF_X1 U1900 ( .A(n474), .Z(n477) );
  BUF_X1 U1901 ( .A(n481), .Z(n478) );
  BUF_X1 U1902 ( .A(n481), .Z(n479) );
  BUF_X1 U1903 ( .A(n481), .Z(n480) );
  INV_X1 U1904 ( .A(n448), .ZN(n481) );
  INV_X1 U1905 ( .A(n4870), .ZN(n482) );
  INV_X1 U1906 ( .A(n4870), .ZN(n483) );
  INV_X1 U1907 ( .A(n4870), .ZN(n484) );
  INV_X1 U1908 ( .A(n4870), .ZN(n485) );
  INV_X1 U1909 ( .A(addr[4]), .ZN(n1540) );
  INV_X1 U1910 ( .A(addr[4]), .ZN(n1541) );
  INV_X1 U1911 ( .A(addr[4]), .ZN(n1542) );
  INV_X1 U1912 ( .A(addr[5]), .ZN(n1563) );
  INV_X1 U1913 ( .A(addr[6]), .ZN(n1575) );
  INV_X1 U1914 ( .A(n1580), .ZN(n1576) );
  INV_X1 U1915 ( .A(n1583), .ZN(n1577) );
endmodule


module gng_smul_16_18_sadd_37_DW01_add_0 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [37:2] carry;

  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .S(SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module gng_smul_16_18_sadd_37_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .A(n70), .ZN(n13) );
  INV_X1 U3 ( .A(n62), .ZN(n11) );
  INV_X1 U4 ( .A(n54), .ZN(n9) );
  INV_X1 U5 ( .A(n46), .ZN(n7) );
  INV_X1 U6 ( .A(n38), .ZN(n5) );
  INV_X1 U7 ( .A(n30), .ZN(n3) );
  INV_X1 U8 ( .A(n32), .ZN(n4) );
  INV_X1 U9 ( .A(n24), .ZN(n2) );
  INV_X1 U10 ( .A(n72), .ZN(n14) );
  INV_X1 U11 ( .A(n64), .ZN(n12) );
  INV_X1 U12 ( .A(n56), .ZN(n10) );
  INV_X1 U13 ( .A(n48), .ZN(n8) );
  INV_X1 U14 ( .A(n40), .ZN(n6) );
  INV_X1 U15 ( .A(n22), .ZN(n1) );
  INV_X1 U16 ( .A(n78), .ZN(n15) );
  INV_X1 U17 ( .A(n80), .ZN(n16) );
  INV_X1 U18 ( .A(n84), .ZN(SUM[14]) );
  XOR2_X1 U19 ( .A(n18), .B(n19), .Z(SUM[31]) );
  AOI21_X1 U20 ( .B1(n20), .B2(n1), .A(n21), .ZN(n19) );
  XNOR2_X1 U21 ( .A(B[31]), .B(A[31]), .ZN(n18) );
  XOR2_X1 U22 ( .A(n20), .B(n23), .Z(SUM[30]) );
  NOR2_X1 U23 ( .A1(n21), .A2(n22), .ZN(n23) );
  NOR2_X1 U24 ( .A1(B[30]), .A2(A[30]), .ZN(n22) );
  AND2_X1 U25 ( .A1(B[30]), .A2(A[30]), .ZN(n21) );
  OAI21_X1 U26 ( .B1(n24), .B2(n25), .A(n26), .ZN(n20) );
  XOR2_X1 U27 ( .A(n27), .B(n25), .Z(SUM[29]) );
  AOI21_X1 U28 ( .B1(n3), .B2(n28), .A(n29), .ZN(n25) );
  NAND2_X1 U29 ( .A1(n2), .A2(n26), .ZN(n27) );
  NAND2_X1 U30 ( .A1(B[29]), .A2(A[29]), .ZN(n26) );
  NOR2_X1 U31 ( .A1(B[29]), .A2(A[29]), .ZN(n24) );
  XOR2_X1 U32 ( .A(n28), .B(n31), .Z(SUM[28]) );
  NOR2_X1 U33 ( .A1(n29), .A2(n30), .ZN(n31) );
  NOR2_X1 U34 ( .A1(B[28]), .A2(A[28]), .ZN(n30) );
  AND2_X1 U35 ( .A1(B[28]), .A2(A[28]), .ZN(n29) );
  OAI21_X1 U36 ( .B1(n32), .B2(n33), .A(n34), .ZN(n28) );
  XOR2_X1 U37 ( .A(n35), .B(n33), .Z(SUM[27]) );
  AOI21_X1 U38 ( .B1(n5), .B2(n36), .A(n37), .ZN(n33) );
  NAND2_X1 U39 ( .A1(n4), .A2(n34), .ZN(n35) );
  NAND2_X1 U40 ( .A1(B[27]), .A2(A[27]), .ZN(n34) );
  NOR2_X1 U41 ( .A1(B[27]), .A2(A[27]), .ZN(n32) );
  XOR2_X1 U42 ( .A(n36), .B(n39), .Z(SUM[26]) );
  NOR2_X1 U43 ( .A1(n37), .A2(n38), .ZN(n39) );
  NOR2_X1 U44 ( .A1(B[26]), .A2(A[26]), .ZN(n38) );
  AND2_X1 U45 ( .A1(B[26]), .A2(A[26]), .ZN(n37) );
  OAI21_X1 U46 ( .B1(n40), .B2(n41), .A(n42), .ZN(n36) );
  XOR2_X1 U47 ( .A(n43), .B(n41), .Z(SUM[25]) );
  AOI21_X1 U48 ( .B1(n7), .B2(n44), .A(n45), .ZN(n41) );
  NAND2_X1 U49 ( .A1(n6), .A2(n42), .ZN(n43) );
  NAND2_X1 U50 ( .A1(B[25]), .A2(A[25]), .ZN(n42) );
  NOR2_X1 U51 ( .A1(B[25]), .A2(A[25]), .ZN(n40) );
  XOR2_X1 U52 ( .A(n44), .B(n47), .Z(SUM[24]) );
  NOR2_X1 U53 ( .A1(n45), .A2(n46), .ZN(n47) );
  NOR2_X1 U54 ( .A1(B[24]), .A2(A[24]), .ZN(n46) );
  AND2_X1 U55 ( .A1(B[24]), .A2(A[24]), .ZN(n45) );
  OAI21_X1 U56 ( .B1(n48), .B2(n49), .A(n50), .ZN(n44) );
  XOR2_X1 U57 ( .A(n51), .B(n49), .Z(SUM[23]) );
  AOI21_X1 U58 ( .B1(n9), .B2(n52), .A(n53), .ZN(n49) );
  NAND2_X1 U59 ( .A1(n8), .A2(n50), .ZN(n51) );
  NAND2_X1 U60 ( .A1(B[23]), .A2(A[23]), .ZN(n50) );
  NOR2_X1 U61 ( .A1(B[23]), .A2(A[23]), .ZN(n48) );
  XOR2_X1 U62 ( .A(n52), .B(n55), .Z(SUM[22]) );
  NOR2_X1 U63 ( .A1(n53), .A2(n54), .ZN(n55) );
  NOR2_X1 U64 ( .A1(B[22]), .A2(A[22]), .ZN(n54) );
  AND2_X1 U65 ( .A1(B[22]), .A2(A[22]), .ZN(n53) );
  OAI21_X1 U66 ( .B1(n56), .B2(n57), .A(n58), .ZN(n52) );
  XOR2_X1 U67 ( .A(n59), .B(n57), .Z(SUM[21]) );
  AOI21_X1 U68 ( .B1(n11), .B2(n60), .A(n61), .ZN(n57) );
  NAND2_X1 U69 ( .A1(n10), .A2(n58), .ZN(n59) );
  NAND2_X1 U70 ( .A1(B[21]), .A2(A[21]), .ZN(n58) );
  NOR2_X1 U71 ( .A1(B[21]), .A2(A[21]), .ZN(n56) );
  XOR2_X1 U72 ( .A(n60), .B(n63), .Z(SUM[20]) );
  NOR2_X1 U73 ( .A1(n61), .A2(n62), .ZN(n63) );
  NOR2_X1 U74 ( .A1(B[20]), .A2(A[20]), .ZN(n62) );
  AND2_X1 U75 ( .A1(B[20]), .A2(A[20]), .ZN(n61) );
  OAI21_X1 U76 ( .B1(n64), .B2(n65), .A(n66), .ZN(n60) );
  XOR2_X1 U77 ( .A(n67), .B(n65), .Z(SUM[19]) );
  AOI21_X1 U78 ( .B1(n13), .B2(n68), .A(n69), .ZN(n65) );
  NAND2_X1 U79 ( .A1(n12), .A2(n66), .ZN(n67) );
  NAND2_X1 U80 ( .A1(B[19]), .A2(A[19]), .ZN(n66) );
  NOR2_X1 U81 ( .A1(B[19]), .A2(A[19]), .ZN(n64) );
  XOR2_X1 U82 ( .A(n68), .B(n71), .Z(SUM[18]) );
  NOR2_X1 U83 ( .A1(n69), .A2(n70), .ZN(n71) );
  NOR2_X1 U84 ( .A1(B[18]), .A2(A[18]), .ZN(n70) );
  AND2_X1 U85 ( .A1(B[18]), .A2(A[18]), .ZN(n69) );
  OAI21_X1 U86 ( .B1(n72), .B2(n73), .A(n74), .ZN(n68) );
  XOR2_X1 U87 ( .A(n75), .B(n73), .Z(SUM[17]) );
  AOI21_X1 U88 ( .B1(n15), .B2(n76), .A(n77), .ZN(n73) );
  NAND2_X1 U89 ( .A1(n14), .A2(n74), .ZN(n75) );
  NAND2_X1 U90 ( .A1(B[17]), .A2(A[17]), .ZN(n74) );
  NOR2_X1 U91 ( .A1(B[17]), .A2(A[17]), .ZN(n72) );
  XOR2_X1 U92 ( .A(n76), .B(n79), .Z(SUM[16]) );
  NOR2_X1 U93 ( .A1(n77), .A2(n78), .ZN(n79) );
  NOR2_X1 U94 ( .A1(B[16]), .A2(A[16]), .ZN(n78) );
  AND2_X1 U95 ( .A1(B[16]), .A2(A[16]), .ZN(n77) );
  OAI21_X1 U96 ( .B1(n80), .B2(n81), .A(n82), .ZN(n76) );
  XOR2_X1 U97 ( .A(n81), .B(n83), .Z(SUM[15]) );
  NAND2_X1 U98 ( .A1(n16), .A2(n82), .ZN(n83) );
  NAND2_X1 U99 ( .A1(B[15]), .A2(A[15]), .ZN(n82) );
  NOR2_X1 U100 ( .A1(B[15]), .A2(A[15]), .ZN(n80) );
  OAI21_X1 U101 ( .B1(B[14]), .B2(A[14]), .A(n81), .ZN(n84) );
  NAND2_X1 U102 ( .A1(B[14]), .A2(A[14]), .ZN(n81) );
endmodule


module gng_smul_16_18_sadd_37_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [17:0] B;
  output [33:0] PRODUCT;
  input TC;
  wire   ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_, ab_15__13_,
         ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_,
         ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_,
         ab_15__0_, ab_14__17_, ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_,
         ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_,
         ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_,
         ab_14__0_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_, ab_13__13_,
         ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_,
         ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_,
         ab_13__0_, ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_,
         ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_,
         ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_,
         ab_11__0_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_, ab_10__13_,
         ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_, ab_10__7_,
         ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_, ab_10__1_,
         ab_10__0_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__17_,
         ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_, ab_7__11_,
         ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_,
         ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__17_, ab_6__16_,
         ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_, ab_6__11_, ab_6__10_,
         ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_,
         ab_6__2_, ab_6__1_, ab_6__0_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_,
         ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_,
         ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_,
         ab_4__0_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_, ab_3__13_,
         ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_, ab_3__7_,
         ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_,
         ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_, ab_2__13_, ab_2__12_,
         ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__17_,
         ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_,
         ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_,
         ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__17_, CARRYB_15__16_, CARRYB_15__15_,
         CARRYB_15__14_, CARRYB_15__13_, CARRYB_15__12_, CARRYB_15__11_,
         CARRYB_15__10_, CARRYB_15__9_, CARRYB_15__8_, CARRYB_15__7_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__16_, CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_,
         CARRYB_13__12_, CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_,
         CARRYB_13__8_, CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_, CARRYB_9__13_,
         CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_, CARRYB_9__9_,
         CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_, CARRYB_9__4_,
         CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__16_,
         CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_, CARRYB_7__12_,
         CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_, CARRYB_7__8_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__16_,
         CARRYB_4__15_, CARRYB_4__14_, CARRYB_4__13_, CARRYB_4__12_,
         CARRYB_4__11_, CARRYB_4__10_, CARRYB_4__9_, CARRYB_4__8_,
         CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_15__0_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__16_, SUMB_13__15_, SUMB_13__14_,
         SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_, SUMB_13__9_,
         SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__16_,
         SUMB_11__15_, SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_,
         SUMB_11__10_, SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_,
         SUMB_11__5_, SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_,
         SUMB_10__16_, SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_,
         SUMB_10__11_, SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__16_, SUMB_8__15_, SUMB_8__14_,
         SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_, SUMB_8__9_,
         SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__16_,
         SUMB_6__15_, SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_,
         SUMB_6__10_, SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_,
         SUMB_6__5_, SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_,
         SUMB_5__16_, SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_,
         SUMB_5__11_, SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__16_, SUMB_3__15_, SUMB_3__14_,
         SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_, SUMB_3__9_,
         SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, A1_15_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_,
         A1_2_, A1_1_, A1_0_, A2_16_, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104;

  FA_X1 S14_17_0 ( .A(B[17]), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(A2_16_), 
        .S(A1_15_) );
  FA_X1 S4_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(SUMB_15__0_) );
  FA_X1 S4_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S4_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S4_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S4_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S4_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S4_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S4_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S4_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S4_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S4_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S4_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S4_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S4_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S4_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S4_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S5_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(ab_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S14_17 ( .A(n71), .B(n87), .CI(ab_15__17_), .CO(CARRYB_15__17_), .S(
        SUMB_15__17_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S3_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(ab_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S3_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(ab_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S3_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(ab_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S3_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(ab_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S3_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(ab_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S3_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(ab_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S3_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(ab_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S3_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(ab_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S3_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(ab_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S3_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(ab_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S3_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(ab_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S3_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(ab_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n17), .CI(n34), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n16), .CI(n33), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n15), .CI(n31), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n14), .CI(n30), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n13), .CI(n29), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n12), .CI(n28), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(n11), .CI(n27), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(n10), .CI(n26), .CO(CARRYB_2__7_), .S(
        SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(n9), .CI(n25), .CO(CARRYB_2__8_), .S(
        SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(n8), .CI(n24), .CO(CARRYB_2__9_), .S(
        SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(n7), .CI(n23), .CO(CARRYB_2__10_), .S(
        SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(n6), .CI(n22), .CO(CARRYB_2__11_), .S(
        SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(n5), .CI(n21), .CO(CARRYB_2__12_), .S(
        SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(n4), .CI(n20), .CO(CARRYB_2__13_), .S(
        SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(n3), .CI(n19), .CO(CARRYB_2__14_), .S(
        SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(n2), .CI(n32), .CO(CARRYB_2__15_), .S(
        SUMB_2__15_) );
  FA_X1 S3_2_16 ( .A(ab_2__16_), .B(n18), .CI(ab_1__17_), .CO(CARRYB_2__16_), 
        .S(SUMB_2__16_) );
  gng_smul_16_18_sadd_37_DW01_add_1 FS_1 ( .A({n70, n48, n67, n47, n66, n46, 
        n65, n45, n64, n44, n63, n43, n62, n37, n42, n36, A1_15_, n38, n69, 
        A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, 
        A1_3_, A1_2_, A1_1_, A1_0_}), .B({n49, n61, n60, n59, n58, n57, n56, 
        n55, n54, n53, n52, n51, n50, n41, n40, A2_16_, n39, n68, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[33:2]) );
  AND2_X1 U2 ( .A1(ab_0__16_), .A2(ab_1__15_), .ZN(n2) );
  AND2_X1 U3 ( .A1(ab_0__15_), .A2(ab_1__14_), .ZN(n3) );
  AND2_X1 U4 ( .A1(ab_0__14_), .A2(ab_1__13_), .ZN(n4) );
  AND2_X1 U5 ( .A1(ab_0__13_), .A2(ab_1__12_), .ZN(n5) );
  AND2_X1 U6 ( .A1(ab_0__12_), .A2(ab_1__11_), .ZN(n6) );
  AND2_X1 U7 ( .A1(ab_0__11_), .A2(ab_1__10_), .ZN(n7) );
  AND2_X1 U8 ( .A1(ab_0__10_), .A2(ab_1__9_), .ZN(n8) );
  AND2_X1 U9 ( .A1(ab_0__9_), .A2(ab_1__8_), .ZN(n9) );
  AND2_X1 U10 ( .A1(ab_0__8_), .A2(ab_1__7_), .ZN(n10) );
  AND2_X1 U11 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n11) );
  AND2_X1 U12 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n12) );
  AND2_X1 U13 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n13) );
  AND2_X1 U14 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n14) );
  AND2_X1 U15 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n15) );
  AND2_X1 U16 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n16) );
  AND2_X1 U17 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n17) );
  AND2_X1 U18 ( .A1(ab_0__17_), .A2(ab_1__16_), .ZN(n18) );
  XOR2_X1 U19 ( .A(ab_1__15_), .B(ab_0__16_), .Z(n19) );
  XOR2_X1 U20 ( .A(ab_1__14_), .B(ab_0__15_), .Z(n20) );
  XOR2_X1 U21 ( .A(ab_1__13_), .B(ab_0__14_), .Z(n21) );
  XOR2_X1 U22 ( .A(ab_1__12_), .B(ab_0__13_), .Z(n22) );
  XOR2_X1 U23 ( .A(ab_1__11_), .B(ab_0__12_), .Z(n23) );
  XOR2_X1 U24 ( .A(ab_1__10_), .B(ab_0__11_), .Z(n24) );
  XOR2_X1 U25 ( .A(ab_1__9_), .B(ab_0__10_), .Z(n25) );
  XOR2_X1 U26 ( .A(ab_1__8_), .B(ab_0__9_), .Z(n26) );
  XOR2_X1 U27 ( .A(ab_1__7_), .B(ab_0__8_), .Z(n27) );
  XOR2_X1 U28 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n28) );
  XOR2_X1 U29 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n29) );
  XOR2_X1 U30 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n30) );
  XOR2_X1 U31 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n31) );
  XOR2_X1 U32 ( .A(ab_1__16_), .B(ab_0__17_), .Z(n32) );
  XOR2_X1 U33 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n33) );
  XOR2_X1 U34 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n34) );
  INV_X1 U35 ( .A(CARRYB_15__17_), .ZN(n70) );
  XOR2_X1 U36 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U37 ( .A(CARRYB_15__2_), .B(SUMB_15__3_), .Z(n36) );
  XOR2_X1 U38 ( .A(CARRYB_15__4_), .B(SUMB_15__5_), .Z(n37) );
  XOR2_X1 U39 ( .A(CARRYB_15__0_), .B(SUMB_15__1_), .Z(n38) );
  AND2_X1 U40 ( .A1(CARRYB_15__0_), .A2(SUMB_15__1_), .ZN(n39) );
  AND2_X1 U41 ( .A1(CARRYB_15__2_), .A2(SUMB_15__3_), .ZN(n40) );
  AND2_X1 U42 ( .A1(CARRYB_15__3_), .A2(SUMB_15__4_), .ZN(n41) );
  XOR2_X1 U43 ( .A(CARRYB_15__3_), .B(SUMB_15__4_), .Z(n42) );
  XOR2_X1 U44 ( .A(CARRYB_15__6_), .B(SUMB_15__7_), .Z(n43) );
  XOR2_X1 U45 ( .A(CARRYB_15__8_), .B(SUMB_15__9_), .Z(n44) );
  XOR2_X1 U46 ( .A(CARRYB_15__10_), .B(SUMB_15__11_), .Z(n45) );
  XOR2_X1 U47 ( .A(CARRYB_15__12_), .B(SUMB_15__13_), .Z(n46) );
  XOR2_X1 U48 ( .A(CARRYB_15__14_), .B(SUMB_15__15_), .Z(n47) );
  XOR2_X1 U49 ( .A(CARRYB_15__16_), .B(SUMB_15__17_), .Z(n48) );
  AND2_X1 U50 ( .A1(CARRYB_15__16_), .A2(SUMB_15__17_), .ZN(n49) );
  AND2_X1 U51 ( .A1(CARRYB_15__4_), .A2(SUMB_15__5_), .ZN(n50) );
  AND2_X1 U52 ( .A1(CARRYB_15__5_), .A2(SUMB_15__6_), .ZN(n51) );
  AND2_X1 U53 ( .A1(CARRYB_15__6_), .A2(SUMB_15__7_), .ZN(n52) );
  AND2_X1 U54 ( .A1(CARRYB_15__7_), .A2(SUMB_15__8_), .ZN(n53) );
  AND2_X1 U55 ( .A1(CARRYB_15__8_), .A2(SUMB_15__9_), .ZN(n54) );
  AND2_X1 U56 ( .A1(CARRYB_15__9_), .A2(SUMB_15__10_), .ZN(n55) );
  AND2_X1 U57 ( .A1(CARRYB_15__10_), .A2(SUMB_15__11_), .ZN(n56) );
  AND2_X1 U58 ( .A1(CARRYB_15__11_), .A2(SUMB_15__12_), .ZN(n57) );
  AND2_X1 U59 ( .A1(CARRYB_15__12_), .A2(SUMB_15__13_), .ZN(n58) );
  AND2_X1 U60 ( .A1(CARRYB_15__13_), .A2(SUMB_15__14_), .ZN(n59) );
  AND2_X1 U61 ( .A1(CARRYB_15__14_), .A2(SUMB_15__15_), .ZN(n60) );
  AND2_X1 U62 ( .A1(CARRYB_15__15_), .A2(SUMB_15__16_), .ZN(n61) );
  XOR2_X1 U63 ( .A(CARRYB_15__5_), .B(SUMB_15__6_), .Z(n62) );
  XOR2_X1 U64 ( .A(CARRYB_15__7_), .B(SUMB_15__8_), .Z(n63) );
  XOR2_X1 U65 ( .A(CARRYB_15__9_), .B(SUMB_15__10_), .Z(n64) );
  XOR2_X1 U66 ( .A(CARRYB_15__11_), .B(SUMB_15__12_), .Z(n65) );
  XOR2_X1 U67 ( .A(CARRYB_15__13_), .B(SUMB_15__14_), .Z(n66) );
  XOR2_X1 U68 ( .A(CARRYB_15__15_), .B(SUMB_15__16_), .Z(n67) );
  INV_X1 U69 ( .A(B[17]), .ZN(n87) );
  INV_X1 U70 ( .A(A[0]), .ZN(n86) );
  INV_X1 U71 ( .A(A[1]), .ZN(n85) );
  INV_X1 U72 ( .A(A[3]), .ZN(n83) );
  INV_X1 U73 ( .A(A[2]), .ZN(n84) );
  INV_X1 U74 ( .A(B[8]), .ZN(n96) );
  INV_X1 U75 ( .A(B[7]), .ZN(n97) );
  INV_X1 U76 ( .A(B[6]), .ZN(n98) );
  INV_X1 U77 ( .A(B[5]), .ZN(n99) );
  INV_X1 U78 ( .A(B[4]), .ZN(n100) );
  INV_X1 U79 ( .A(B[3]), .ZN(n101) );
  INV_X1 U80 ( .A(B[2]), .ZN(n102) );
  INV_X1 U81 ( .A(B[10]), .ZN(n94) );
  INV_X1 U82 ( .A(B[9]), .ZN(n95) );
  INV_X1 U83 ( .A(B[12]), .ZN(n92) );
  INV_X1 U84 ( .A(B[11]), .ZN(n93) );
  INV_X1 U85 ( .A(B[14]), .ZN(n90) );
  INV_X1 U86 ( .A(B[13]), .ZN(n91) );
  INV_X1 U87 ( .A(B[16]), .ZN(n88) );
  INV_X1 U88 ( .A(B[15]), .ZN(n89) );
  AND2_X1 U89 ( .A1(A[15]), .A2(SUMB_15__0_), .ZN(n68) );
  INV_X1 U90 ( .A(A[9]), .ZN(n77) );
  INV_X1 U91 ( .A(A[4]), .ZN(n82) );
  INV_X1 U92 ( .A(A[5]), .ZN(n81) );
  INV_X1 U93 ( .A(A[6]), .ZN(n80) );
  INV_X1 U94 ( .A(A[7]), .ZN(n79) );
  INV_X1 U95 ( .A(A[8]), .ZN(n78) );
  INV_X1 U96 ( .A(A[10]), .ZN(n76) );
  INV_X1 U97 ( .A(A[11]), .ZN(n75) );
  INV_X1 U98 ( .A(A[12]), .ZN(n74) );
  INV_X1 U99 ( .A(B[1]), .ZN(n103) );
  INV_X1 U100 ( .A(B[0]), .ZN(n104) );
  XOR2_X1 U101 ( .A(A[15]), .B(SUMB_15__0_), .Z(n69) );
  INV_X1 U102 ( .A(A[15]), .ZN(n71) );
  INV_X1 U103 ( .A(A[13]), .ZN(n73) );
  INV_X1 U104 ( .A(A[14]), .ZN(n72) );
  NOR2_X1 U105 ( .A1(n77), .A2(n95), .ZN(ab_9__9_) );
  NOR2_X1 U106 ( .A1(n77), .A2(n96), .ZN(ab_9__8_) );
  NOR2_X1 U107 ( .A1(n77), .A2(n97), .ZN(ab_9__7_) );
  NOR2_X1 U108 ( .A1(n77), .A2(n98), .ZN(ab_9__6_) );
  NOR2_X1 U109 ( .A1(n77), .A2(n99), .ZN(ab_9__5_) );
  NOR2_X1 U110 ( .A1(n77), .A2(n100), .ZN(ab_9__4_) );
  NOR2_X1 U111 ( .A1(n77), .A2(n101), .ZN(ab_9__3_) );
  NOR2_X1 U112 ( .A1(n77), .A2(n102), .ZN(ab_9__2_) );
  NOR2_X1 U113 ( .A1(n77), .A2(n103), .ZN(ab_9__1_) );
  NOR2_X1 U114 ( .A1(A[9]), .A2(n87), .ZN(ab_9__17_) );
  NOR2_X1 U115 ( .A1(n77), .A2(n88), .ZN(ab_9__16_) );
  NOR2_X1 U116 ( .A1(n77), .A2(n89), .ZN(ab_9__15_) );
  NOR2_X1 U117 ( .A1(n77), .A2(n90), .ZN(ab_9__14_) );
  NOR2_X1 U118 ( .A1(n77), .A2(n91), .ZN(ab_9__13_) );
  NOR2_X1 U119 ( .A1(n77), .A2(n92), .ZN(ab_9__12_) );
  NOR2_X1 U120 ( .A1(n77), .A2(n93), .ZN(ab_9__11_) );
  NOR2_X1 U121 ( .A1(n77), .A2(n94), .ZN(ab_9__10_) );
  NOR2_X1 U122 ( .A1(n77), .A2(n104), .ZN(ab_9__0_) );
  NOR2_X1 U123 ( .A1(n95), .A2(n78), .ZN(ab_8__9_) );
  NOR2_X1 U124 ( .A1(n96), .A2(n78), .ZN(ab_8__8_) );
  NOR2_X1 U125 ( .A1(n97), .A2(n78), .ZN(ab_8__7_) );
  NOR2_X1 U126 ( .A1(n98), .A2(n78), .ZN(ab_8__6_) );
  NOR2_X1 U127 ( .A1(n99), .A2(n78), .ZN(ab_8__5_) );
  NOR2_X1 U128 ( .A1(n100), .A2(n78), .ZN(ab_8__4_) );
  NOR2_X1 U129 ( .A1(n101), .A2(n78), .ZN(ab_8__3_) );
  NOR2_X1 U130 ( .A1(n102), .A2(n78), .ZN(ab_8__2_) );
  NOR2_X1 U131 ( .A1(n103), .A2(n78), .ZN(ab_8__1_) );
  NOR2_X1 U132 ( .A1(A[8]), .A2(n87), .ZN(ab_8__17_) );
  NOR2_X1 U133 ( .A1(n88), .A2(n78), .ZN(ab_8__16_) );
  NOR2_X1 U134 ( .A1(n89), .A2(n78), .ZN(ab_8__15_) );
  NOR2_X1 U135 ( .A1(n90), .A2(n78), .ZN(ab_8__14_) );
  NOR2_X1 U136 ( .A1(n91), .A2(n78), .ZN(ab_8__13_) );
  NOR2_X1 U137 ( .A1(n92), .A2(n78), .ZN(ab_8__12_) );
  NOR2_X1 U138 ( .A1(n93), .A2(n78), .ZN(ab_8__11_) );
  NOR2_X1 U139 ( .A1(n94), .A2(n78), .ZN(ab_8__10_) );
  NOR2_X1 U140 ( .A1(n104), .A2(n78), .ZN(ab_8__0_) );
  NOR2_X1 U141 ( .A1(n95), .A2(n79), .ZN(ab_7__9_) );
  NOR2_X1 U142 ( .A1(n96), .A2(n79), .ZN(ab_7__8_) );
  NOR2_X1 U143 ( .A1(n97), .A2(n79), .ZN(ab_7__7_) );
  NOR2_X1 U144 ( .A1(n98), .A2(n79), .ZN(ab_7__6_) );
  NOR2_X1 U145 ( .A1(n99), .A2(n79), .ZN(ab_7__5_) );
  NOR2_X1 U146 ( .A1(n100), .A2(n79), .ZN(ab_7__4_) );
  NOR2_X1 U147 ( .A1(n101), .A2(n79), .ZN(ab_7__3_) );
  NOR2_X1 U148 ( .A1(n102), .A2(n79), .ZN(ab_7__2_) );
  NOR2_X1 U149 ( .A1(n103), .A2(n79), .ZN(ab_7__1_) );
  NOR2_X1 U150 ( .A1(A[7]), .A2(n87), .ZN(ab_7__17_) );
  NOR2_X1 U151 ( .A1(n88), .A2(n79), .ZN(ab_7__16_) );
  NOR2_X1 U152 ( .A1(n89), .A2(n79), .ZN(ab_7__15_) );
  NOR2_X1 U153 ( .A1(n90), .A2(n79), .ZN(ab_7__14_) );
  NOR2_X1 U154 ( .A1(n91), .A2(n79), .ZN(ab_7__13_) );
  NOR2_X1 U155 ( .A1(n92), .A2(n79), .ZN(ab_7__12_) );
  NOR2_X1 U156 ( .A1(n93), .A2(n79), .ZN(ab_7__11_) );
  NOR2_X1 U157 ( .A1(n94), .A2(n79), .ZN(ab_7__10_) );
  NOR2_X1 U158 ( .A1(n104), .A2(n79), .ZN(ab_7__0_) );
  NOR2_X1 U159 ( .A1(n95), .A2(n80), .ZN(ab_6__9_) );
  NOR2_X1 U160 ( .A1(n96), .A2(n80), .ZN(ab_6__8_) );
  NOR2_X1 U161 ( .A1(n97), .A2(n80), .ZN(ab_6__7_) );
  NOR2_X1 U162 ( .A1(n98), .A2(n80), .ZN(ab_6__6_) );
  NOR2_X1 U163 ( .A1(n99), .A2(n80), .ZN(ab_6__5_) );
  NOR2_X1 U164 ( .A1(n100), .A2(n80), .ZN(ab_6__4_) );
  NOR2_X1 U165 ( .A1(n101), .A2(n80), .ZN(ab_6__3_) );
  NOR2_X1 U166 ( .A1(n102), .A2(n80), .ZN(ab_6__2_) );
  NOR2_X1 U167 ( .A1(n103), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U168 ( .A1(A[6]), .A2(n87), .ZN(ab_6__17_) );
  NOR2_X1 U169 ( .A1(n88), .A2(n80), .ZN(ab_6__16_) );
  NOR2_X1 U170 ( .A1(n89), .A2(n80), .ZN(ab_6__15_) );
  NOR2_X1 U171 ( .A1(n90), .A2(n80), .ZN(ab_6__14_) );
  NOR2_X1 U172 ( .A1(n91), .A2(n80), .ZN(ab_6__13_) );
  NOR2_X1 U173 ( .A1(n92), .A2(n80), .ZN(ab_6__12_) );
  NOR2_X1 U174 ( .A1(n93), .A2(n80), .ZN(ab_6__11_) );
  NOR2_X1 U175 ( .A1(n94), .A2(n80), .ZN(ab_6__10_) );
  NOR2_X1 U176 ( .A1(n104), .A2(n80), .ZN(ab_6__0_) );
  NOR2_X1 U177 ( .A1(n95), .A2(n81), .ZN(ab_5__9_) );
  NOR2_X1 U178 ( .A1(n96), .A2(n81), .ZN(ab_5__8_) );
  NOR2_X1 U179 ( .A1(n97), .A2(n81), .ZN(ab_5__7_) );
  NOR2_X1 U180 ( .A1(n98), .A2(n81), .ZN(ab_5__6_) );
  NOR2_X1 U181 ( .A1(n99), .A2(n81), .ZN(ab_5__5_) );
  NOR2_X1 U182 ( .A1(n100), .A2(n81), .ZN(ab_5__4_) );
  NOR2_X1 U183 ( .A1(n101), .A2(n81), .ZN(ab_5__3_) );
  NOR2_X1 U184 ( .A1(n102), .A2(n81), .ZN(ab_5__2_) );
  NOR2_X1 U185 ( .A1(n103), .A2(n81), .ZN(ab_5__1_) );
  NOR2_X1 U186 ( .A1(A[5]), .A2(n87), .ZN(ab_5__17_) );
  NOR2_X1 U187 ( .A1(n88), .A2(n81), .ZN(ab_5__16_) );
  NOR2_X1 U188 ( .A1(n89), .A2(n81), .ZN(ab_5__15_) );
  NOR2_X1 U189 ( .A1(n90), .A2(n81), .ZN(ab_5__14_) );
  NOR2_X1 U190 ( .A1(n91), .A2(n81), .ZN(ab_5__13_) );
  NOR2_X1 U191 ( .A1(n92), .A2(n81), .ZN(ab_5__12_) );
  NOR2_X1 U192 ( .A1(n93), .A2(n81), .ZN(ab_5__11_) );
  NOR2_X1 U193 ( .A1(n94), .A2(n81), .ZN(ab_5__10_) );
  NOR2_X1 U194 ( .A1(n104), .A2(n81), .ZN(ab_5__0_) );
  NOR2_X1 U195 ( .A1(n95), .A2(n82), .ZN(ab_4__9_) );
  NOR2_X1 U196 ( .A1(n96), .A2(n82), .ZN(ab_4__8_) );
  NOR2_X1 U197 ( .A1(n97), .A2(n82), .ZN(ab_4__7_) );
  NOR2_X1 U198 ( .A1(n98), .A2(n82), .ZN(ab_4__6_) );
  NOR2_X1 U199 ( .A1(n99), .A2(n82), .ZN(ab_4__5_) );
  NOR2_X1 U200 ( .A1(n100), .A2(n82), .ZN(ab_4__4_) );
  NOR2_X1 U201 ( .A1(n101), .A2(n82), .ZN(ab_4__3_) );
  NOR2_X1 U202 ( .A1(n102), .A2(n82), .ZN(ab_4__2_) );
  NOR2_X1 U203 ( .A1(n103), .A2(n82), .ZN(ab_4__1_) );
  NOR2_X1 U204 ( .A1(A[4]), .A2(n87), .ZN(ab_4__17_) );
  NOR2_X1 U205 ( .A1(n88), .A2(n82), .ZN(ab_4__16_) );
  NOR2_X1 U206 ( .A1(n89), .A2(n82), .ZN(ab_4__15_) );
  NOR2_X1 U207 ( .A1(n90), .A2(n82), .ZN(ab_4__14_) );
  NOR2_X1 U208 ( .A1(n91), .A2(n82), .ZN(ab_4__13_) );
  NOR2_X1 U209 ( .A1(n92), .A2(n82), .ZN(ab_4__12_) );
  NOR2_X1 U210 ( .A1(n93), .A2(n82), .ZN(ab_4__11_) );
  NOR2_X1 U211 ( .A1(n94), .A2(n82), .ZN(ab_4__10_) );
  NOR2_X1 U212 ( .A1(n104), .A2(n82), .ZN(ab_4__0_) );
  NOR2_X1 U213 ( .A1(n95), .A2(n83), .ZN(ab_3__9_) );
  NOR2_X1 U214 ( .A1(n96), .A2(n83), .ZN(ab_3__8_) );
  NOR2_X1 U215 ( .A1(n97), .A2(n83), .ZN(ab_3__7_) );
  NOR2_X1 U216 ( .A1(n98), .A2(n83), .ZN(ab_3__6_) );
  NOR2_X1 U217 ( .A1(n99), .A2(n83), .ZN(ab_3__5_) );
  NOR2_X1 U218 ( .A1(n100), .A2(n83), .ZN(ab_3__4_) );
  NOR2_X1 U219 ( .A1(n101), .A2(n83), .ZN(ab_3__3_) );
  NOR2_X1 U220 ( .A1(n102), .A2(n83), .ZN(ab_3__2_) );
  NOR2_X1 U221 ( .A1(n103), .A2(n83), .ZN(ab_3__1_) );
  NOR2_X1 U222 ( .A1(A[3]), .A2(n87), .ZN(ab_3__17_) );
  NOR2_X1 U223 ( .A1(n88), .A2(n83), .ZN(ab_3__16_) );
  NOR2_X1 U224 ( .A1(n89), .A2(n83), .ZN(ab_3__15_) );
  NOR2_X1 U225 ( .A1(n90), .A2(n83), .ZN(ab_3__14_) );
  NOR2_X1 U226 ( .A1(n91), .A2(n83), .ZN(ab_3__13_) );
  NOR2_X1 U227 ( .A1(n92), .A2(n83), .ZN(ab_3__12_) );
  NOR2_X1 U228 ( .A1(n93), .A2(n83), .ZN(ab_3__11_) );
  NOR2_X1 U229 ( .A1(n94), .A2(n83), .ZN(ab_3__10_) );
  NOR2_X1 U230 ( .A1(n104), .A2(n83), .ZN(ab_3__0_) );
  NOR2_X1 U231 ( .A1(n95), .A2(n84), .ZN(ab_2__9_) );
  NOR2_X1 U232 ( .A1(n96), .A2(n84), .ZN(ab_2__8_) );
  NOR2_X1 U233 ( .A1(n97), .A2(n84), .ZN(ab_2__7_) );
  NOR2_X1 U234 ( .A1(n98), .A2(n84), .ZN(ab_2__6_) );
  NOR2_X1 U235 ( .A1(n99), .A2(n84), .ZN(ab_2__5_) );
  NOR2_X1 U236 ( .A1(n100), .A2(n84), .ZN(ab_2__4_) );
  NOR2_X1 U237 ( .A1(n101), .A2(n84), .ZN(ab_2__3_) );
  NOR2_X1 U238 ( .A1(n102), .A2(n84), .ZN(ab_2__2_) );
  NOR2_X1 U239 ( .A1(n103), .A2(n84), .ZN(ab_2__1_) );
  NOR2_X1 U240 ( .A1(A[2]), .A2(n87), .ZN(ab_2__17_) );
  NOR2_X1 U241 ( .A1(n88), .A2(n84), .ZN(ab_2__16_) );
  NOR2_X1 U242 ( .A1(n89), .A2(n84), .ZN(ab_2__15_) );
  NOR2_X1 U243 ( .A1(n90), .A2(n84), .ZN(ab_2__14_) );
  NOR2_X1 U244 ( .A1(n91), .A2(n84), .ZN(ab_2__13_) );
  NOR2_X1 U245 ( .A1(n92), .A2(n84), .ZN(ab_2__12_) );
  NOR2_X1 U246 ( .A1(n93), .A2(n84), .ZN(ab_2__11_) );
  NOR2_X1 U247 ( .A1(n94), .A2(n84), .ZN(ab_2__10_) );
  NOR2_X1 U248 ( .A1(n104), .A2(n84), .ZN(ab_2__0_) );
  NOR2_X1 U249 ( .A1(n95), .A2(n85), .ZN(ab_1__9_) );
  NOR2_X1 U250 ( .A1(n96), .A2(n85), .ZN(ab_1__8_) );
  NOR2_X1 U251 ( .A1(n97), .A2(n85), .ZN(ab_1__7_) );
  NOR2_X1 U252 ( .A1(n98), .A2(n85), .ZN(ab_1__6_) );
  NOR2_X1 U253 ( .A1(n99), .A2(n85), .ZN(ab_1__5_) );
  NOR2_X1 U254 ( .A1(n100), .A2(n85), .ZN(ab_1__4_) );
  NOR2_X1 U255 ( .A1(n101), .A2(n85), .ZN(ab_1__3_) );
  NOR2_X1 U256 ( .A1(n102), .A2(n85), .ZN(ab_1__2_) );
  NOR2_X1 U257 ( .A1(n103), .A2(n85), .ZN(ab_1__1_) );
  NOR2_X1 U258 ( .A1(A[1]), .A2(n87), .ZN(ab_1__17_) );
  NOR2_X1 U259 ( .A1(n88), .A2(n85), .ZN(ab_1__16_) );
  NOR2_X1 U260 ( .A1(n89), .A2(n85), .ZN(ab_1__15_) );
  NOR2_X1 U261 ( .A1(n90), .A2(n85), .ZN(ab_1__14_) );
  NOR2_X1 U262 ( .A1(n91), .A2(n85), .ZN(ab_1__13_) );
  NOR2_X1 U263 ( .A1(n92), .A2(n85), .ZN(ab_1__12_) );
  NOR2_X1 U264 ( .A1(n93), .A2(n85), .ZN(ab_1__11_) );
  NOR2_X1 U265 ( .A1(n94), .A2(n85), .ZN(ab_1__10_) );
  NOR2_X1 U266 ( .A1(n104), .A2(n85), .ZN(ab_1__0_) );
  NOR2_X1 U267 ( .A1(B[9]), .A2(n71), .ZN(ab_15__9_) );
  NOR2_X1 U268 ( .A1(B[8]), .A2(n71), .ZN(ab_15__8_) );
  NOR2_X1 U269 ( .A1(B[7]), .A2(n71), .ZN(ab_15__7_) );
  NOR2_X1 U270 ( .A1(B[6]), .A2(n71), .ZN(ab_15__6_) );
  NOR2_X1 U271 ( .A1(B[5]), .A2(n71), .ZN(ab_15__5_) );
  NOR2_X1 U272 ( .A1(B[4]), .A2(n71), .ZN(ab_15__4_) );
  NOR2_X1 U273 ( .A1(B[3]), .A2(n71), .ZN(ab_15__3_) );
  NOR2_X1 U274 ( .A1(B[2]), .A2(n71), .ZN(ab_15__2_) );
  NOR2_X1 U275 ( .A1(B[1]), .A2(n71), .ZN(ab_15__1_) );
  NOR2_X1 U276 ( .A1(n87), .A2(n71), .ZN(ab_15__17_) );
  NOR2_X1 U277 ( .A1(B[16]), .A2(n71), .ZN(ab_15__16_) );
  NOR2_X1 U278 ( .A1(B[15]), .A2(n71), .ZN(ab_15__15_) );
  NOR2_X1 U279 ( .A1(B[14]), .A2(n71), .ZN(ab_15__14_) );
  NOR2_X1 U280 ( .A1(B[13]), .A2(n71), .ZN(ab_15__13_) );
  NOR2_X1 U281 ( .A1(B[12]), .A2(n71), .ZN(ab_15__12_) );
  NOR2_X1 U282 ( .A1(B[11]), .A2(n71), .ZN(ab_15__11_) );
  NOR2_X1 U283 ( .A1(B[10]), .A2(n71), .ZN(ab_15__10_) );
  NOR2_X1 U284 ( .A1(B[0]), .A2(n71), .ZN(ab_15__0_) );
  NOR2_X1 U285 ( .A1(n95), .A2(n72), .ZN(ab_14__9_) );
  NOR2_X1 U286 ( .A1(n96), .A2(n72), .ZN(ab_14__8_) );
  NOR2_X1 U287 ( .A1(n97), .A2(n72), .ZN(ab_14__7_) );
  NOR2_X1 U288 ( .A1(n98), .A2(n72), .ZN(ab_14__6_) );
  NOR2_X1 U289 ( .A1(n99), .A2(n72), .ZN(ab_14__5_) );
  NOR2_X1 U290 ( .A1(n100), .A2(n72), .ZN(ab_14__4_) );
  NOR2_X1 U291 ( .A1(n101), .A2(n72), .ZN(ab_14__3_) );
  NOR2_X1 U292 ( .A1(n102), .A2(n72), .ZN(ab_14__2_) );
  NOR2_X1 U293 ( .A1(n103), .A2(n72), .ZN(ab_14__1_) );
  NOR2_X1 U294 ( .A1(A[14]), .A2(n87), .ZN(ab_14__17_) );
  NOR2_X1 U295 ( .A1(n88), .A2(n72), .ZN(ab_14__16_) );
  NOR2_X1 U296 ( .A1(n89), .A2(n72), .ZN(ab_14__15_) );
  NOR2_X1 U297 ( .A1(n90), .A2(n72), .ZN(ab_14__14_) );
  NOR2_X1 U298 ( .A1(n91), .A2(n72), .ZN(ab_14__13_) );
  NOR2_X1 U299 ( .A1(n92), .A2(n72), .ZN(ab_14__12_) );
  NOR2_X1 U300 ( .A1(n93), .A2(n72), .ZN(ab_14__11_) );
  NOR2_X1 U301 ( .A1(n94), .A2(n72), .ZN(ab_14__10_) );
  NOR2_X1 U302 ( .A1(n104), .A2(n72), .ZN(ab_14__0_) );
  NOR2_X1 U303 ( .A1(n95), .A2(n73), .ZN(ab_13__9_) );
  NOR2_X1 U304 ( .A1(n96), .A2(n73), .ZN(ab_13__8_) );
  NOR2_X1 U305 ( .A1(n97), .A2(n73), .ZN(ab_13__7_) );
  NOR2_X1 U306 ( .A1(n98), .A2(n73), .ZN(ab_13__6_) );
  NOR2_X1 U307 ( .A1(n99), .A2(n73), .ZN(ab_13__5_) );
  NOR2_X1 U308 ( .A1(n100), .A2(n73), .ZN(ab_13__4_) );
  NOR2_X1 U309 ( .A1(n101), .A2(n73), .ZN(ab_13__3_) );
  NOR2_X1 U310 ( .A1(n102), .A2(n73), .ZN(ab_13__2_) );
  NOR2_X1 U311 ( .A1(n103), .A2(n73), .ZN(ab_13__1_) );
  NOR2_X1 U312 ( .A1(A[13]), .A2(n87), .ZN(ab_13__17_) );
  NOR2_X1 U313 ( .A1(n88), .A2(n73), .ZN(ab_13__16_) );
  NOR2_X1 U314 ( .A1(n89), .A2(n73), .ZN(ab_13__15_) );
  NOR2_X1 U315 ( .A1(n90), .A2(n73), .ZN(ab_13__14_) );
  NOR2_X1 U316 ( .A1(n91), .A2(n73), .ZN(ab_13__13_) );
  NOR2_X1 U317 ( .A1(n92), .A2(n73), .ZN(ab_13__12_) );
  NOR2_X1 U318 ( .A1(n93), .A2(n73), .ZN(ab_13__11_) );
  NOR2_X1 U319 ( .A1(n94), .A2(n73), .ZN(ab_13__10_) );
  NOR2_X1 U320 ( .A1(n104), .A2(n73), .ZN(ab_13__0_) );
  NOR2_X1 U321 ( .A1(n95), .A2(n74), .ZN(ab_12__9_) );
  NOR2_X1 U322 ( .A1(n96), .A2(n74), .ZN(ab_12__8_) );
  NOR2_X1 U323 ( .A1(n97), .A2(n74), .ZN(ab_12__7_) );
  NOR2_X1 U324 ( .A1(n98), .A2(n74), .ZN(ab_12__6_) );
  NOR2_X1 U325 ( .A1(n99), .A2(n74), .ZN(ab_12__5_) );
  NOR2_X1 U326 ( .A1(n100), .A2(n74), .ZN(ab_12__4_) );
  NOR2_X1 U327 ( .A1(n101), .A2(n74), .ZN(ab_12__3_) );
  NOR2_X1 U328 ( .A1(n102), .A2(n74), .ZN(ab_12__2_) );
  NOR2_X1 U329 ( .A1(n103), .A2(n74), .ZN(ab_12__1_) );
  NOR2_X1 U330 ( .A1(A[12]), .A2(n87), .ZN(ab_12__17_) );
  NOR2_X1 U331 ( .A1(n88), .A2(n74), .ZN(ab_12__16_) );
  NOR2_X1 U332 ( .A1(n89), .A2(n74), .ZN(ab_12__15_) );
  NOR2_X1 U333 ( .A1(n90), .A2(n74), .ZN(ab_12__14_) );
  NOR2_X1 U334 ( .A1(n91), .A2(n74), .ZN(ab_12__13_) );
  NOR2_X1 U335 ( .A1(n92), .A2(n74), .ZN(ab_12__12_) );
  NOR2_X1 U336 ( .A1(n93), .A2(n74), .ZN(ab_12__11_) );
  NOR2_X1 U337 ( .A1(n94), .A2(n74), .ZN(ab_12__10_) );
  NOR2_X1 U338 ( .A1(n104), .A2(n74), .ZN(ab_12__0_) );
  NOR2_X1 U339 ( .A1(n95), .A2(n75), .ZN(ab_11__9_) );
  NOR2_X1 U340 ( .A1(n96), .A2(n75), .ZN(ab_11__8_) );
  NOR2_X1 U341 ( .A1(n97), .A2(n75), .ZN(ab_11__7_) );
  NOR2_X1 U342 ( .A1(n98), .A2(n75), .ZN(ab_11__6_) );
  NOR2_X1 U343 ( .A1(n99), .A2(n75), .ZN(ab_11__5_) );
  NOR2_X1 U344 ( .A1(n100), .A2(n75), .ZN(ab_11__4_) );
  NOR2_X1 U345 ( .A1(n101), .A2(n75), .ZN(ab_11__3_) );
  NOR2_X1 U346 ( .A1(n102), .A2(n75), .ZN(ab_11__2_) );
  NOR2_X1 U347 ( .A1(n103), .A2(n75), .ZN(ab_11__1_) );
  NOR2_X1 U348 ( .A1(A[11]), .A2(n87), .ZN(ab_11__17_) );
  NOR2_X1 U349 ( .A1(n88), .A2(n75), .ZN(ab_11__16_) );
  NOR2_X1 U350 ( .A1(n89), .A2(n75), .ZN(ab_11__15_) );
  NOR2_X1 U351 ( .A1(n90), .A2(n75), .ZN(ab_11__14_) );
  NOR2_X1 U352 ( .A1(n91), .A2(n75), .ZN(ab_11__13_) );
  NOR2_X1 U353 ( .A1(n92), .A2(n75), .ZN(ab_11__12_) );
  NOR2_X1 U354 ( .A1(n93), .A2(n75), .ZN(ab_11__11_) );
  NOR2_X1 U355 ( .A1(n94), .A2(n75), .ZN(ab_11__10_) );
  NOR2_X1 U356 ( .A1(n104), .A2(n75), .ZN(ab_11__0_) );
  NOR2_X1 U357 ( .A1(n95), .A2(n76), .ZN(ab_10__9_) );
  NOR2_X1 U358 ( .A1(n96), .A2(n76), .ZN(ab_10__8_) );
  NOR2_X1 U359 ( .A1(n97), .A2(n76), .ZN(ab_10__7_) );
  NOR2_X1 U360 ( .A1(n98), .A2(n76), .ZN(ab_10__6_) );
  NOR2_X1 U361 ( .A1(n99), .A2(n76), .ZN(ab_10__5_) );
  NOR2_X1 U362 ( .A1(n100), .A2(n76), .ZN(ab_10__4_) );
  NOR2_X1 U363 ( .A1(n101), .A2(n76), .ZN(ab_10__3_) );
  NOR2_X1 U364 ( .A1(n102), .A2(n76), .ZN(ab_10__2_) );
  NOR2_X1 U365 ( .A1(n103), .A2(n76), .ZN(ab_10__1_) );
  NOR2_X1 U366 ( .A1(A[10]), .A2(n87), .ZN(ab_10__17_) );
  NOR2_X1 U367 ( .A1(n88), .A2(n76), .ZN(ab_10__16_) );
  NOR2_X1 U368 ( .A1(n89), .A2(n76), .ZN(ab_10__15_) );
  NOR2_X1 U369 ( .A1(n90), .A2(n76), .ZN(ab_10__14_) );
  NOR2_X1 U370 ( .A1(n91), .A2(n76), .ZN(ab_10__13_) );
  NOR2_X1 U371 ( .A1(n92), .A2(n76), .ZN(ab_10__12_) );
  NOR2_X1 U372 ( .A1(n93), .A2(n76), .ZN(ab_10__11_) );
  NOR2_X1 U373 ( .A1(n94), .A2(n76), .ZN(ab_10__10_) );
  NOR2_X1 U374 ( .A1(n104), .A2(n76), .ZN(ab_10__0_) );
  NOR2_X1 U375 ( .A1(n95), .A2(n86), .ZN(ab_0__9_) );
  NOR2_X1 U376 ( .A1(n96), .A2(n86), .ZN(ab_0__8_) );
  NOR2_X1 U377 ( .A1(n97), .A2(n86), .ZN(ab_0__7_) );
  NOR2_X1 U378 ( .A1(n98), .A2(n86), .ZN(ab_0__6_) );
  NOR2_X1 U379 ( .A1(n99), .A2(n86), .ZN(ab_0__5_) );
  NOR2_X1 U380 ( .A1(n100), .A2(n86), .ZN(ab_0__4_) );
  NOR2_X1 U381 ( .A1(n101), .A2(n86), .ZN(ab_0__3_) );
  NOR2_X1 U382 ( .A1(n102), .A2(n86), .ZN(ab_0__2_) );
  NOR2_X1 U383 ( .A1(n103), .A2(n86), .ZN(ab_0__1_) );
  NOR2_X1 U384 ( .A1(A[0]), .A2(n87), .ZN(ab_0__17_) );
  NOR2_X1 U385 ( .A1(n88), .A2(n86), .ZN(ab_0__16_) );
  NOR2_X1 U386 ( .A1(n89), .A2(n86), .ZN(ab_0__15_) );
  NOR2_X1 U387 ( .A1(n90), .A2(n86), .ZN(ab_0__14_) );
  NOR2_X1 U388 ( .A1(n91), .A2(n86), .ZN(ab_0__13_) );
  NOR2_X1 U389 ( .A1(n92), .A2(n86), .ZN(ab_0__12_) );
  NOR2_X1 U390 ( .A1(n93), .A2(n86), .ZN(ab_0__11_) );
  NOR2_X1 U391 ( .A1(n94), .A2(n86), .ZN(ab_0__10_) );
  NOR2_X1 U392 ( .A1(n104), .A2(n86), .ZN(PRODUCT[0]) );
endmodule


module gng_smul_16_18_sadd_37 ( clk, a, b, c, p );
  input [15:0] a;
  input [17:0] b;
  input [36:0] c;
  output [37:0] p;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33;
  wire   [15:0] a_reg;
  wire   [17:0] b_reg;
  wire   [36:0] c_reg;
  wire   [33:0] prod;
  wire   [37:0] sum;

  DFF_X1 a_reg_reg_15_ ( .D(a[15]), .CK(clk), .Q(a_reg[15]) );
  DFF_X1 a_reg_reg_14_ ( .D(a[14]), .CK(clk), .Q(a_reg[14]) );
  DFF_X1 a_reg_reg_13_ ( .D(a[13]), .CK(clk), .Q(a_reg[13]) );
  DFF_X1 a_reg_reg_12_ ( .D(a[12]), .CK(clk), .Q(a_reg[12]) );
  DFF_X1 a_reg_reg_11_ ( .D(a[11]), .CK(clk), .Q(a_reg[11]) );
  DFF_X1 a_reg_reg_10_ ( .D(a[10]), .CK(clk), .Q(a_reg[10]) );
  DFF_X1 a_reg_reg_9_ ( .D(a[9]), .CK(clk), .Q(a_reg[9]) );
  DFF_X1 a_reg_reg_8_ ( .D(a[8]), .CK(clk), .Q(a_reg[8]) );
  DFF_X1 a_reg_reg_7_ ( .D(a[7]), .CK(clk), .Q(a_reg[7]) );
  DFF_X1 a_reg_reg_6_ ( .D(a[6]), .CK(clk), .Q(a_reg[6]) );
  DFF_X1 a_reg_reg_5_ ( .D(a[5]), .CK(clk), .Q(a_reg[5]) );
  DFF_X1 a_reg_reg_4_ ( .D(a[4]), .CK(clk), .Q(a_reg[4]) );
  DFF_X1 a_reg_reg_3_ ( .D(a[3]), .CK(clk), .Q(a_reg[3]) );
  DFF_X1 a_reg_reg_2_ ( .D(a[2]), .CK(clk), .Q(a_reg[2]) );
  DFF_X1 a_reg_reg_1_ ( .D(a[1]), .CK(clk), .Q(a_reg[1]) );
  DFF_X1 a_reg_reg_0_ ( .D(a[0]), .CK(clk), .Q(a_reg[0]) );
  DFF_X1 b_reg_reg_17_ ( .D(b[17]), .CK(clk), .Q(b_reg[17]) );
  DFF_X1 b_reg_reg_16_ ( .D(b[16]), .CK(clk), .Q(b_reg[16]) );
  DFF_X1 b_reg_reg_15_ ( .D(b[15]), .CK(clk), .Q(b_reg[15]) );
  DFF_X1 b_reg_reg_14_ ( .D(b[14]), .CK(clk), .Q(b_reg[14]) );
  DFF_X1 b_reg_reg_13_ ( .D(b[13]), .CK(clk), .Q(b_reg[13]) );
  DFF_X1 b_reg_reg_12_ ( .D(b[12]), .CK(clk), .Q(b_reg[12]) );
  DFF_X1 b_reg_reg_11_ ( .D(b[11]), .CK(clk), .Q(b_reg[11]) );
  DFF_X1 b_reg_reg_10_ ( .D(b[10]), .CK(clk), .Q(b_reg[10]) );
  DFF_X1 b_reg_reg_9_ ( .D(b[9]), .CK(clk), .Q(b_reg[9]) );
  DFF_X1 b_reg_reg_8_ ( .D(b[8]), .CK(clk), .Q(b_reg[8]) );
  DFF_X1 b_reg_reg_7_ ( .D(b[7]), .CK(clk), .Q(b_reg[7]) );
  DFF_X1 b_reg_reg_6_ ( .D(b[6]), .CK(clk), .Q(b_reg[6]) );
  DFF_X1 b_reg_reg_5_ ( .D(b[5]), .CK(clk), .Q(b_reg[5]) );
  DFF_X1 b_reg_reg_4_ ( .D(b[4]), .CK(clk), .Q(b_reg[4]) );
  DFF_X1 b_reg_reg_3_ ( .D(b[3]), .CK(clk), .Q(b_reg[3]) );
  DFF_X1 b_reg_reg_2_ ( .D(b[2]), .CK(clk), .Q(b_reg[2]) );
  DFF_X1 b_reg_reg_1_ ( .D(b[1]), .CK(clk), .Q(b_reg[1]) );
  DFF_X1 b_reg_reg_0_ ( .D(b[0]), .CK(clk), .Q(b_reg[0]) );
  DFF_X1 c_reg_reg_36_ ( .D(c[36]), .CK(clk), .Q(c_reg[36]) );
  DFF_X1 c_reg_reg_35_ ( .D(c[35]), .CK(clk), .Q(c_reg[35]) );
  DFF_X1 c_reg_reg_34_ ( .D(c[34]), .CK(clk), .Q(c_reg[34]) );
  DFF_X1 c_reg_reg_33_ ( .D(c[33]), .CK(clk), .Q(c_reg[33]) );
  DFF_X1 c_reg_reg_32_ ( .D(c[32]), .CK(clk), .Q(c_reg[32]) );
  DFF_X1 c_reg_reg_31_ ( .D(c[31]), .CK(clk), .Q(c_reg[31]) );
  DFF_X1 c_reg_reg_30_ ( .D(c[30]), .CK(clk), .Q(c_reg[30]) );
  DFF_X1 c_reg_reg_29_ ( .D(c[29]), .CK(clk), .Q(c_reg[29]) );
  DFF_X1 c_reg_reg_28_ ( .D(c[28]), .CK(clk), .Q(c_reg[28]) );
  DFF_X1 c_reg_reg_27_ ( .D(c[27]), .CK(clk), .Q(c_reg[27]) );
  DFF_X1 c_reg_reg_26_ ( .D(c[26]), .CK(clk), .Q(c_reg[26]) );
  DFF_X1 c_reg_reg_25_ ( .D(c[25]), .CK(clk), .Q(c_reg[25]) );
  DFF_X1 c_reg_reg_24_ ( .D(c[24]), .CK(clk), .Q(c_reg[24]) );
  DFF_X1 c_reg_reg_23_ ( .D(c[23]), .CK(clk), .Q(c_reg[23]) );
  DFF_X1 c_reg_reg_22_ ( .D(c[22]), .CK(clk), .Q(c_reg[22]) );
  DFF_X1 c_reg_reg_21_ ( .D(c[21]), .CK(clk), .Q(c_reg[21]) );
  DFF_X1 c_reg_reg_20_ ( .D(c[20]), .CK(clk), .Q(c_reg[20]) );
  DFF_X1 c_reg_reg_19_ ( .D(c[19]), .CK(clk), .Q(c_reg[19]) );
  DFF_X1 c_reg_reg_18_ ( .D(c[18]), .CK(clk), .Q(c_reg[18]) );
  DFF_X1 c_reg_reg_17_ ( .D(c[17]), .CK(clk), .Q(c_reg[17]) );
  DFF_X1 c_reg_reg_16_ ( .D(c[16]), .CK(clk), .Q(c_reg[16]) );
  DFF_X1 c_reg_reg_15_ ( .D(c[15]), .CK(clk), .Q(c_reg[15]) );
  DFF_X1 c_reg_reg_14_ ( .D(c[14]), .CK(clk), .Q(c_reg[14]) );
  DFF_X1 c_reg_reg_13_ ( .D(c[13]), .CK(clk), .Q(c_reg[13]) );
  DFF_X1 c_reg_reg_12_ ( .D(c[12]), .CK(clk), .Q(c_reg[12]) );
  DFF_X1 c_reg_reg_11_ ( .D(c[11]), .CK(clk), .Q(c_reg[11]) );
  DFF_X1 c_reg_reg_10_ ( .D(c[10]), .CK(clk), .Q(c_reg[10]) );
  DFF_X1 c_reg_reg_9_ ( .D(c[9]), .CK(clk), .Q(c_reg[9]) );
  DFF_X1 c_reg_reg_8_ ( .D(c[8]), .CK(clk), .Q(c_reg[8]) );
  DFF_X1 c_reg_reg_7_ ( .D(c[7]), .CK(clk), .Q(c_reg[7]) );
  DFF_X1 c_reg_reg_6_ ( .D(c[6]), .CK(clk), .Q(c_reg[6]) );
  DFF_X1 c_reg_reg_5_ ( .D(c[5]), .CK(clk), .Q(c_reg[5]) );
  DFF_X1 c_reg_reg_4_ ( .D(c[4]), .CK(clk), .Q(c_reg[4]) );
  DFF_X1 c_reg_reg_3_ ( .D(c[3]), .CK(clk), .Q(c_reg[3]) );
  DFF_X1 c_reg_reg_2_ ( .D(c[2]), .CK(clk), .Q(c_reg[2]) );
  DFF_X1 c_reg_reg_1_ ( .D(c[1]), .CK(clk), .Q(c_reg[1]) );
  DFF_X1 c_reg_reg_0_ ( .D(c[0]), .CK(clk), .Q(c_reg[0]) );
  DFF_X1 prod_reg_33_ ( .D(N33), .CK(clk), .Q(prod[33]) );
  DFF_X1 prod_reg_32_ ( .D(N32), .CK(clk), .Q(prod[32]) );
  DFF_X1 prod_reg_31_ ( .D(N31), .CK(clk), .Q(prod[31]) );
  DFF_X1 prod_reg_30_ ( .D(N30), .CK(clk), .Q(prod[30]) );
  DFF_X1 prod_reg_29_ ( .D(N29), .CK(clk), .Q(prod[29]) );
  DFF_X1 prod_reg_28_ ( .D(N28), .CK(clk), .Q(prod[28]) );
  DFF_X1 prod_reg_27_ ( .D(N27), .CK(clk), .Q(prod[27]) );
  DFF_X1 prod_reg_26_ ( .D(N26), .CK(clk), .Q(prod[26]) );
  DFF_X1 prod_reg_25_ ( .D(N25), .CK(clk), .Q(prod[25]) );
  DFF_X1 prod_reg_24_ ( .D(N24), .CK(clk), .Q(prod[24]) );
  DFF_X1 prod_reg_23_ ( .D(N23), .CK(clk), .Q(prod[23]) );
  DFF_X1 prod_reg_22_ ( .D(N22), .CK(clk), .Q(prod[22]) );
  DFF_X1 prod_reg_21_ ( .D(N21), .CK(clk), .Q(prod[21]) );
  DFF_X1 prod_reg_20_ ( .D(N20), .CK(clk), .Q(prod[20]) );
  DFF_X1 prod_reg_19_ ( .D(N19), .CK(clk), .Q(prod[19]) );
  DFF_X1 prod_reg_18_ ( .D(N18), .CK(clk), .Q(prod[18]) );
  DFF_X1 prod_reg_17_ ( .D(N17), .CK(clk), .Q(prod[17]) );
  DFF_X1 prod_reg_16_ ( .D(N16), .CK(clk), .Q(prod[16]) );
  DFF_X1 prod_reg_15_ ( .D(N15), .CK(clk), .Q(prod[15]) );
  DFF_X1 prod_reg_14_ ( .D(N14), .CK(clk), .Q(prod[14]) );
  DFF_X1 prod_reg_13_ ( .D(N13), .CK(clk), .Q(prod[13]) );
  DFF_X1 prod_reg_12_ ( .D(N12), .CK(clk), .Q(prod[12]) );
  DFF_X1 prod_reg_11_ ( .D(N11), .CK(clk), .Q(prod[11]) );
  DFF_X1 prod_reg_10_ ( .D(N10), .CK(clk), .Q(prod[10]) );
  DFF_X1 prod_reg_9_ ( .D(N9), .CK(clk), .Q(prod[9]) );
  DFF_X1 prod_reg_8_ ( .D(N8), .CK(clk), .Q(prod[8]) );
  DFF_X1 prod_reg_7_ ( .D(N7), .CK(clk), .Q(prod[7]) );
  DFF_X1 prod_reg_6_ ( .D(N6), .CK(clk), .Q(prod[6]) );
  DFF_X1 prod_reg_5_ ( .D(N5), .CK(clk), .Q(prod[5]) );
  DFF_X1 prod_reg_4_ ( .D(N4), .CK(clk), .Q(prod[4]) );
  DFF_X1 prod_reg_3_ ( .D(N3), .CK(clk), .Q(prod[3]) );
  DFF_X1 prod_reg_2_ ( .D(N2), .CK(clk), .Q(prod[2]) );
  DFF_X1 prod_reg_1_ ( .D(N1), .CK(clk), .Q(prod[1]) );
  DFF_X1 prod_reg_0_ ( .D(N0), .CK(clk), .Q(prod[0]) );
  DFF_X1 result_reg_37_ ( .D(sum[37]), .CK(clk), .Q(p[37]) );
  DFF_X1 result_reg_36_ ( .D(sum[36]), .CK(clk), .Q(p[36]) );
  DFF_X1 result_reg_35_ ( .D(sum[35]), .CK(clk), .Q(p[35]) );
  DFF_X1 result_reg_34_ ( .D(sum[34]), .CK(clk), .Q(p[34]) );
  DFF_X1 result_reg_33_ ( .D(sum[33]), .CK(clk), .Q(p[33]) );
  DFF_X1 result_reg_32_ ( .D(sum[32]), .CK(clk), .Q(p[32]) );
  DFF_X1 result_reg_31_ ( .D(sum[31]), .CK(clk), .Q(p[31]) );
  DFF_X1 result_reg_30_ ( .D(sum[30]), .CK(clk), .Q(p[30]) );
  DFF_X1 result_reg_29_ ( .D(sum[29]), .CK(clk), .Q(p[29]) );
  DFF_X1 result_reg_28_ ( .D(sum[28]), .CK(clk), .Q(p[28]) );
  DFF_X1 result_reg_27_ ( .D(sum[27]), .CK(clk), .Q(p[27]) );
  DFF_X1 result_reg_26_ ( .D(sum[26]), .CK(clk), .Q(p[26]) );
  DFF_X1 result_reg_25_ ( .D(sum[25]), .CK(clk), .Q(p[25]) );
  DFF_X1 result_reg_24_ ( .D(sum[24]), .CK(clk), .Q(p[24]) );
  DFF_X1 result_reg_23_ ( .D(sum[23]), .CK(clk), .Q(p[23]) );
  DFF_X1 result_reg_22_ ( .D(sum[22]), .CK(clk), .Q(p[22]) );
  DFF_X1 result_reg_21_ ( .D(sum[21]), .CK(clk), .Q(p[21]) );
  DFF_X1 result_reg_20_ ( .D(sum[20]), .CK(clk), .Q(p[20]) );
  DFF_X1 result_reg_19_ ( .D(sum[19]), .CK(clk), .Q(p[19]) );
  DFF_X1 result_reg_18_ ( .D(sum[18]), .CK(clk), .Q(p[18]) );
  DFF_X1 result_reg_17_ ( .D(sum[17]), .CK(clk), .Q(p[17]) );
  DFF_X1 result_reg_16_ ( .D(sum[16]), .CK(clk), .Q(p[16]) );
  DFF_X1 result_reg_15_ ( .D(sum[15]), .CK(clk), .Q(p[15]) );
  DFF_X1 result_reg_14_ ( .D(sum[14]), .CK(clk), .Q(p[14]) );
  DFF_X1 result_reg_13_ ( .D(sum[13]), .CK(clk), .Q(p[13]) );
  DFF_X1 result_reg_12_ ( .D(sum[12]), .CK(clk), .Q(p[12]) );
  DFF_X1 result_reg_11_ ( .D(sum[11]), .CK(clk), .Q(p[11]) );
  DFF_X1 result_reg_10_ ( .D(sum[10]), .CK(clk), .Q(p[10]) );
  DFF_X1 result_reg_9_ ( .D(sum[9]), .CK(clk), .Q(p[9]) );
  DFF_X1 result_reg_8_ ( .D(sum[8]), .CK(clk), .Q(p[8]) );
  DFF_X1 result_reg_7_ ( .D(sum[7]), .CK(clk), .Q(p[7]) );
  DFF_X1 result_reg_6_ ( .D(sum[6]), .CK(clk), .Q(p[6]) );
  DFF_X1 result_reg_5_ ( .D(sum[5]), .CK(clk), .Q(p[5]) );
  DFF_X1 result_reg_4_ ( .D(sum[4]), .CK(clk), .Q(p[4]) );
  DFF_X1 result_reg_3_ ( .D(sum[3]), .CK(clk), .Q(p[3]) );
  DFF_X1 result_reg_2_ ( .D(sum[2]), .CK(clk), .Q(p[2]) );
  DFF_X1 result_reg_1_ ( .D(sum[1]), .CK(clk), .Q(p[1]) );
  DFF_X1 result_reg_0_ ( .D(sum[0]), .CK(clk), .Q(p[0]) );
  gng_smul_16_18_sadd_37_DW01_add_0 add_69 ( .A({c_reg[36], c_reg}), .B({
        prod[33], prod[33], prod[33], prod[33], prod}), .CI(1'b0), .SUM(sum)
         );
  gng_smul_16_18_sadd_37_DW02_mult_0 mult_66 ( .A(a_reg), .B(b_reg), .TC(1'b1), 
        .PRODUCT({N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4, N3, N2, N1, N0}) );
endmodule


module gng_smul_16_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .A(n70), .ZN(n13) );
  INV_X1 U3 ( .A(n62), .ZN(n11) );
  INV_X1 U4 ( .A(n54), .ZN(n9) );
  INV_X1 U5 ( .A(n46), .ZN(n7) );
  INV_X1 U6 ( .A(n38), .ZN(n5) );
  INV_X1 U7 ( .A(n30), .ZN(n3) );
  INV_X1 U8 ( .A(n32), .ZN(n4) );
  INV_X1 U9 ( .A(n24), .ZN(n2) );
  INV_X1 U10 ( .A(n72), .ZN(n14) );
  INV_X1 U11 ( .A(n64), .ZN(n12) );
  INV_X1 U12 ( .A(n56), .ZN(n10) );
  INV_X1 U13 ( .A(n48), .ZN(n8) );
  INV_X1 U14 ( .A(n40), .ZN(n6) );
  INV_X1 U15 ( .A(n22), .ZN(n1) );
  INV_X1 U16 ( .A(n78), .ZN(n15) );
  INV_X1 U17 ( .A(n80), .ZN(n16) );
  INV_X1 U18 ( .A(n84), .ZN(SUM[14]) );
  XOR2_X1 U19 ( .A(n18), .B(n19), .Z(SUM[31]) );
  AOI21_X1 U20 ( .B1(n20), .B2(n1), .A(n21), .ZN(n19) );
  XNOR2_X1 U21 ( .A(B[31]), .B(A[31]), .ZN(n18) );
  XOR2_X1 U22 ( .A(n20), .B(n23), .Z(SUM[30]) );
  NOR2_X1 U23 ( .A1(n21), .A2(n22), .ZN(n23) );
  NOR2_X1 U24 ( .A1(B[30]), .A2(A[30]), .ZN(n22) );
  AND2_X1 U25 ( .A1(B[30]), .A2(A[30]), .ZN(n21) );
  OAI21_X1 U26 ( .B1(n24), .B2(n25), .A(n26), .ZN(n20) );
  XOR2_X1 U27 ( .A(n27), .B(n25), .Z(SUM[29]) );
  AOI21_X1 U28 ( .B1(n3), .B2(n28), .A(n29), .ZN(n25) );
  NAND2_X1 U29 ( .A1(n2), .A2(n26), .ZN(n27) );
  NAND2_X1 U30 ( .A1(B[29]), .A2(A[29]), .ZN(n26) );
  NOR2_X1 U31 ( .A1(B[29]), .A2(A[29]), .ZN(n24) );
  XOR2_X1 U32 ( .A(n28), .B(n31), .Z(SUM[28]) );
  NOR2_X1 U33 ( .A1(n29), .A2(n30), .ZN(n31) );
  NOR2_X1 U34 ( .A1(B[28]), .A2(A[28]), .ZN(n30) );
  AND2_X1 U35 ( .A1(B[28]), .A2(A[28]), .ZN(n29) );
  OAI21_X1 U36 ( .B1(n32), .B2(n33), .A(n34), .ZN(n28) );
  XOR2_X1 U37 ( .A(n35), .B(n33), .Z(SUM[27]) );
  AOI21_X1 U38 ( .B1(n5), .B2(n36), .A(n37), .ZN(n33) );
  NAND2_X1 U39 ( .A1(n4), .A2(n34), .ZN(n35) );
  NAND2_X1 U40 ( .A1(B[27]), .A2(A[27]), .ZN(n34) );
  NOR2_X1 U41 ( .A1(B[27]), .A2(A[27]), .ZN(n32) );
  XOR2_X1 U42 ( .A(n36), .B(n39), .Z(SUM[26]) );
  NOR2_X1 U43 ( .A1(n37), .A2(n38), .ZN(n39) );
  NOR2_X1 U44 ( .A1(B[26]), .A2(A[26]), .ZN(n38) );
  AND2_X1 U45 ( .A1(B[26]), .A2(A[26]), .ZN(n37) );
  OAI21_X1 U46 ( .B1(n40), .B2(n41), .A(n42), .ZN(n36) );
  XOR2_X1 U47 ( .A(n43), .B(n41), .Z(SUM[25]) );
  AOI21_X1 U48 ( .B1(n7), .B2(n44), .A(n45), .ZN(n41) );
  NAND2_X1 U49 ( .A1(n6), .A2(n42), .ZN(n43) );
  NAND2_X1 U50 ( .A1(B[25]), .A2(A[25]), .ZN(n42) );
  NOR2_X1 U51 ( .A1(B[25]), .A2(A[25]), .ZN(n40) );
  XOR2_X1 U52 ( .A(n44), .B(n47), .Z(SUM[24]) );
  NOR2_X1 U53 ( .A1(n45), .A2(n46), .ZN(n47) );
  NOR2_X1 U54 ( .A1(B[24]), .A2(A[24]), .ZN(n46) );
  AND2_X1 U55 ( .A1(B[24]), .A2(A[24]), .ZN(n45) );
  OAI21_X1 U56 ( .B1(n48), .B2(n49), .A(n50), .ZN(n44) );
  XOR2_X1 U57 ( .A(n51), .B(n49), .Z(SUM[23]) );
  AOI21_X1 U58 ( .B1(n9), .B2(n52), .A(n53), .ZN(n49) );
  NAND2_X1 U59 ( .A1(n8), .A2(n50), .ZN(n51) );
  NAND2_X1 U60 ( .A1(B[23]), .A2(A[23]), .ZN(n50) );
  NOR2_X1 U61 ( .A1(B[23]), .A2(A[23]), .ZN(n48) );
  XOR2_X1 U62 ( .A(n52), .B(n55), .Z(SUM[22]) );
  NOR2_X1 U63 ( .A1(n53), .A2(n54), .ZN(n55) );
  NOR2_X1 U64 ( .A1(B[22]), .A2(A[22]), .ZN(n54) );
  AND2_X1 U65 ( .A1(B[22]), .A2(A[22]), .ZN(n53) );
  OAI21_X1 U66 ( .B1(n56), .B2(n57), .A(n58), .ZN(n52) );
  XOR2_X1 U67 ( .A(n59), .B(n57), .Z(SUM[21]) );
  AOI21_X1 U68 ( .B1(n11), .B2(n60), .A(n61), .ZN(n57) );
  NAND2_X1 U69 ( .A1(n10), .A2(n58), .ZN(n59) );
  NAND2_X1 U70 ( .A1(B[21]), .A2(A[21]), .ZN(n58) );
  NOR2_X1 U71 ( .A1(B[21]), .A2(A[21]), .ZN(n56) );
  XOR2_X1 U72 ( .A(n60), .B(n63), .Z(SUM[20]) );
  NOR2_X1 U73 ( .A1(n61), .A2(n62), .ZN(n63) );
  NOR2_X1 U74 ( .A1(B[20]), .A2(A[20]), .ZN(n62) );
  AND2_X1 U75 ( .A1(B[20]), .A2(A[20]), .ZN(n61) );
  OAI21_X1 U76 ( .B1(n64), .B2(n65), .A(n66), .ZN(n60) );
  XOR2_X1 U77 ( .A(n67), .B(n65), .Z(SUM[19]) );
  AOI21_X1 U78 ( .B1(n13), .B2(n68), .A(n69), .ZN(n65) );
  NAND2_X1 U79 ( .A1(n12), .A2(n66), .ZN(n67) );
  NAND2_X1 U80 ( .A1(B[19]), .A2(A[19]), .ZN(n66) );
  NOR2_X1 U81 ( .A1(B[19]), .A2(A[19]), .ZN(n64) );
  XOR2_X1 U82 ( .A(n68), .B(n71), .Z(SUM[18]) );
  NOR2_X1 U83 ( .A1(n69), .A2(n70), .ZN(n71) );
  NOR2_X1 U84 ( .A1(B[18]), .A2(A[18]), .ZN(n70) );
  AND2_X1 U85 ( .A1(B[18]), .A2(A[18]), .ZN(n69) );
  OAI21_X1 U86 ( .B1(n72), .B2(n73), .A(n74), .ZN(n68) );
  XOR2_X1 U87 ( .A(n75), .B(n73), .Z(SUM[17]) );
  AOI21_X1 U88 ( .B1(n15), .B2(n76), .A(n77), .ZN(n73) );
  NAND2_X1 U89 ( .A1(n14), .A2(n74), .ZN(n75) );
  NAND2_X1 U90 ( .A1(B[17]), .A2(A[17]), .ZN(n74) );
  NOR2_X1 U91 ( .A1(B[17]), .A2(A[17]), .ZN(n72) );
  XOR2_X1 U92 ( .A(n76), .B(n79), .Z(SUM[16]) );
  NOR2_X1 U93 ( .A1(n77), .A2(n78), .ZN(n79) );
  NOR2_X1 U94 ( .A1(B[16]), .A2(A[16]), .ZN(n78) );
  AND2_X1 U95 ( .A1(B[16]), .A2(A[16]), .ZN(n77) );
  OAI21_X1 U96 ( .B1(n80), .B2(n81), .A(n82), .ZN(n76) );
  XOR2_X1 U97 ( .A(n81), .B(n83), .Z(SUM[15]) );
  NAND2_X1 U98 ( .A1(n16), .A2(n82), .ZN(n83) );
  NAND2_X1 U99 ( .A1(B[15]), .A2(A[15]), .ZN(n82) );
  NOR2_X1 U100 ( .A1(B[15]), .A2(A[15]), .ZN(n80) );
  OAI21_X1 U101 ( .B1(B[14]), .B2(A[14]), .A(n81), .ZN(n84) );
  NAND2_X1 U102 ( .A1(B[14]), .A2(A[14]), .ZN(n81) );
endmodule


module gng_smul_16_18_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [17:0] B;
  output [33:0] PRODUCT;
  input TC;
  wire   ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_, ab_15__13_,
         ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_,
         ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_,
         ab_15__0_, ab_14__17_, ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_,
         ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_,
         ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_,
         ab_14__0_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_, ab_13__13_,
         ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_,
         ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_,
         ab_13__0_, ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_,
         ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_,
         ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_,
         ab_11__0_, ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_, ab_10__13_,
         ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_, ab_10__7_,
         ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_, ab_10__1_,
         ab_10__0_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_,
         ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__17_,
         ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_, ab_7__11_,
         ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_,
         ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__17_, ab_6__16_,
         ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_, ab_6__11_, ab_6__10_,
         ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_,
         ab_6__2_, ab_6__1_, ab_6__0_, ab_5__17_, ab_5__16_, ab_5__15_,
         ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_,
         ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_,
         ab_5__1_, ab_5__0_, ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_,
         ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_,
         ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_,
         ab_4__0_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_, ab_3__13_,
         ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_, ab_3__7_,
         ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_,
         ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_, ab_2__13_, ab_2__12_,
         ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__17_,
         ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_,
         ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_,
         ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_, ab_0__17_, ab_0__16_,
         ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_,
         ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_,
         ab_0__2_, ab_0__1_, CARRYB_15__17_, CARRYB_15__16_, CARRYB_15__15_,
         CARRYB_15__14_, CARRYB_15__13_, CARRYB_15__12_, CARRYB_15__11_,
         CARRYB_15__10_, CARRYB_15__9_, CARRYB_15__8_, CARRYB_15__7_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__16_, CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_,
         CARRYB_13__12_, CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_,
         CARRYB_13__8_, CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_, CARRYB_9__13_,
         CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_, CARRYB_9__9_,
         CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_, CARRYB_9__4_,
         CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__16_,
         CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_, CARRYB_7__12_,
         CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_, CARRYB_7__8_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__16_,
         CARRYB_4__15_, CARRYB_4__14_, CARRYB_4__13_, CARRYB_4__12_,
         CARRYB_4__11_, CARRYB_4__10_, CARRYB_4__9_, CARRYB_4__8_,
         CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_15__0_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__16_, SUMB_13__15_, SUMB_13__14_,
         SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_, SUMB_13__9_,
         SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__16_,
         SUMB_11__15_, SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_,
         SUMB_11__10_, SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_,
         SUMB_11__5_, SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_,
         SUMB_10__16_, SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_,
         SUMB_10__11_, SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__16_, SUMB_8__15_, SUMB_8__14_,
         SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_, SUMB_8__9_,
         SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__16_,
         SUMB_6__15_, SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_,
         SUMB_6__10_, SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_,
         SUMB_6__5_, SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_,
         SUMB_5__16_, SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_,
         SUMB_5__11_, SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__16_, SUMB_3__15_, SUMB_3__14_,
         SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_, SUMB_3__9_,
         SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, A1_15_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_,
         A1_2_, A1_1_, A1_0_, A2_16_, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104;

  FA_X1 S14_17_0 ( .A(B[17]), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(A2_16_), 
        .S(A1_15_) );
  FA_X1 S4_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(SUMB_15__0_) );
  FA_X1 S4_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S4_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S4_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S4_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S4_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S4_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S4_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S4_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S4_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S4_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S4_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S4_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S4_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S4_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S4_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S5_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(ab_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S14_17 ( .A(n71), .B(n87), .CI(ab_15__17_), .CO(CARRYB_15__17_), .S(
        SUMB_15__17_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S3_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(ab_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S3_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(ab_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S3_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(ab_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S3_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(ab_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S3_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(ab_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S3_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(ab_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S3_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(ab_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S3_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(ab_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S3_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(ab_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S3_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(ab_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S3_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(ab_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S3_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(ab_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n17), .CI(n34), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n16), .CI(n33), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n15), .CI(n31), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n14), .CI(n30), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n13), .CI(n29), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n12), .CI(n28), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(n11), .CI(n27), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(n10), .CI(n26), .CO(CARRYB_2__7_), .S(
        SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(n9), .CI(n25), .CO(CARRYB_2__8_), .S(
        SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(n8), .CI(n24), .CO(CARRYB_2__9_), .S(
        SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(n7), .CI(n23), .CO(CARRYB_2__10_), .S(
        SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(n6), .CI(n22), .CO(CARRYB_2__11_), .S(
        SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(n5), .CI(n21), .CO(CARRYB_2__12_), .S(
        SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(n4), .CI(n20), .CO(CARRYB_2__13_), .S(
        SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(n3), .CI(n19), .CO(CARRYB_2__14_), .S(
        SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(n2), .CI(n32), .CO(CARRYB_2__15_), .S(
        SUMB_2__15_) );
  FA_X1 S3_2_16 ( .A(ab_2__16_), .B(n18), .CI(ab_1__17_), .CO(CARRYB_2__16_), 
        .S(SUMB_2__16_) );
  gng_smul_16_18_DW01_add_0 FS_1 ( .A({n70, n48, n67, n47, n66, n46, n65, n45, 
        n64, n44, n63, n43, n62, n37, n42, n36, A1_15_, n38, n69, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, 
        A1_1_, A1_0_}), .B({n49, n61, n60, n59, n58, n57, n56, n55, n54, n53, 
        n52, n51, n50, n41, n40, A2_16_, n39, n68, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[33:2]) );
  AND2_X1 U2 ( .A1(ab_0__16_), .A2(ab_1__15_), .ZN(n2) );
  AND2_X1 U3 ( .A1(ab_0__15_), .A2(ab_1__14_), .ZN(n3) );
  AND2_X1 U4 ( .A1(ab_0__14_), .A2(ab_1__13_), .ZN(n4) );
  AND2_X1 U5 ( .A1(ab_0__13_), .A2(ab_1__12_), .ZN(n5) );
  AND2_X1 U6 ( .A1(ab_0__12_), .A2(ab_1__11_), .ZN(n6) );
  AND2_X1 U7 ( .A1(ab_0__11_), .A2(ab_1__10_), .ZN(n7) );
  AND2_X1 U8 ( .A1(ab_0__10_), .A2(ab_1__9_), .ZN(n8) );
  AND2_X1 U9 ( .A1(ab_0__9_), .A2(ab_1__8_), .ZN(n9) );
  AND2_X1 U10 ( .A1(ab_0__8_), .A2(ab_1__7_), .ZN(n10) );
  AND2_X1 U11 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n11) );
  AND2_X1 U12 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n12) );
  AND2_X1 U13 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n13) );
  AND2_X1 U14 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n14) );
  AND2_X1 U15 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n15) );
  AND2_X1 U16 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n16) );
  AND2_X1 U17 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n17) );
  AND2_X1 U18 ( .A1(ab_0__17_), .A2(ab_1__16_), .ZN(n18) );
  XOR2_X1 U19 ( .A(ab_1__15_), .B(ab_0__16_), .Z(n19) );
  XOR2_X1 U20 ( .A(ab_1__14_), .B(ab_0__15_), .Z(n20) );
  XOR2_X1 U21 ( .A(ab_1__13_), .B(ab_0__14_), .Z(n21) );
  XOR2_X1 U22 ( .A(ab_1__12_), .B(ab_0__13_), .Z(n22) );
  XOR2_X1 U23 ( .A(ab_1__11_), .B(ab_0__12_), .Z(n23) );
  XOR2_X1 U24 ( .A(ab_1__10_), .B(ab_0__11_), .Z(n24) );
  XOR2_X1 U25 ( .A(ab_1__9_), .B(ab_0__10_), .Z(n25) );
  XOR2_X1 U26 ( .A(ab_1__8_), .B(ab_0__9_), .Z(n26) );
  XOR2_X1 U27 ( .A(ab_1__7_), .B(ab_0__8_), .Z(n27) );
  XOR2_X1 U28 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n28) );
  XOR2_X1 U29 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n29) );
  XOR2_X1 U30 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n30) );
  XOR2_X1 U31 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n31) );
  XOR2_X1 U32 ( .A(ab_1__16_), .B(ab_0__17_), .Z(n32) );
  XOR2_X1 U33 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n33) );
  XOR2_X1 U34 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n34) );
  INV_X1 U35 ( .A(CARRYB_15__17_), .ZN(n70) );
  XOR2_X1 U36 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U37 ( .A(CARRYB_15__2_), .B(SUMB_15__3_), .Z(n36) );
  XOR2_X1 U38 ( .A(CARRYB_15__4_), .B(SUMB_15__5_), .Z(n37) );
  XOR2_X1 U39 ( .A(CARRYB_15__0_), .B(SUMB_15__1_), .Z(n38) );
  AND2_X1 U40 ( .A1(CARRYB_15__0_), .A2(SUMB_15__1_), .ZN(n39) );
  AND2_X1 U41 ( .A1(CARRYB_15__2_), .A2(SUMB_15__3_), .ZN(n40) );
  AND2_X1 U42 ( .A1(CARRYB_15__3_), .A2(SUMB_15__4_), .ZN(n41) );
  XOR2_X1 U43 ( .A(CARRYB_15__3_), .B(SUMB_15__4_), .Z(n42) );
  XOR2_X1 U44 ( .A(CARRYB_15__6_), .B(SUMB_15__7_), .Z(n43) );
  XOR2_X1 U45 ( .A(CARRYB_15__8_), .B(SUMB_15__9_), .Z(n44) );
  XOR2_X1 U46 ( .A(CARRYB_15__10_), .B(SUMB_15__11_), .Z(n45) );
  XOR2_X1 U47 ( .A(CARRYB_15__12_), .B(SUMB_15__13_), .Z(n46) );
  XOR2_X1 U48 ( .A(CARRYB_15__14_), .B(SUMB_15__15_), .Z(n47) );
  XOR2_X1 U49 ( .A(CARRYB_15__16_), .B(SUMB_15__17_), .Z(n48) );
  AND2_X1 U50 ( .A1(CARRYB_15__16_), .A2(SUMB_15__17_), .ZN(n49) );
  AND2_X1 U51 ( .A1(CARRYB_15__4_), .A2(SUMB_15__5_), .ZN(n50) );
  AND2_X1 U52 ( .A1(CARRYB_15__5_), .A2(SUMB_15__6_), .ZN(n51) );
  AND2_X1 U53 ( .A1(CARRYB_15__6_), .A2(SUMB_15__7_), .ZN(n52) );
  AND2_X1 U54 ( .A1(CARRYB_15__7_), .A2(SUMB_15__8_), .ZN(n53) );
  AND2_X1 U55 ( .A1(CARRYB_15__8_), .A2(SUMB_15__9_), .ZN(n54) );
  AND2_X1 U56 ( .A1(CARRYB_15__9_), .A2(SUMB_15__10_), .ZN(n55) );
  AND2_X1 U57 ( .A1(CARRYB_15__10_), .A2(SUMB_15__11_), .ZN(n56) );
  AND2_X1 U58 ( .A1(CARRYB_15__11_), .A2(SUMB_15__12_), .ZN(n57) );
  AND2_X1 U59 ( .A1(CARRYB_15__12_), .A2(SUMB_15__13_), .ZN(n58) );
  AND2_X1 U60 ( .A1(CARRYB_15__13_), .A2(SUMB_15__14_), .ZN(n59) );
  AND2_X1 U61 ( .A1(CARRYB_15__14_), .A2(SUMB_15__15_), .ZN(n60) );
  AND2_X1 U62 ( .A1(CARRYB_15__15_), .A2(SUMB_15__16_), .ZN(n61) );
  XOR2_X1 U63 ( .A(CARRYB_15__5_), .B(SUMB_15__6_), .Z(n62) );
  XOR2_X1 U64 ( .A(CARRYB_15__7_), .B(SUMB_15__8_), .Z(n63) );
  XOR2_X1 U65 ( .A(CARRYB_15__9_), .B(SUMB_15__10_), .Z(n64) );
  XOR2_X1 U66 ( .A(CARRYB_15__11_), .B(SUMB_15__12_), .Z(n65) );
  XOR2_X1 U67 ( .A(CARRYB_15__13_), .B(SUMB_15__14_), .Z(n66) );
  XOR2_X1 U68 ( .A(CARRYB_15__15_), .B(SUMB_15__16_), .Z(n67) );
  INV_X1 U69 ( .A(B[17]), .ZN(n87) );
  INV_X1 U70 ( .A(A[0]), .ZN(n86) );
  INV_X1 U71 ( .A(A[1]), .ZN(n85) );
  INV_X1 U72 ( .A(A[3]), .ZN(n83) );
  INV_X1 U73 ( .A(A[2]), .ZN(n84) );
  INV_X1 U74 ( .A(B[8]), .ZN(n96) );
  INV_X1 U75 ( .A(B[7]), .ZN(n97) );
  INV_X1 U76 ( .A(B[6]), .ZN(n98) );
  INV_X1 U77 ( .A(B[5]), .ZN(n99) );
  INV_X1 U78 ( .A(B[4]), .ZN(n100) );
  INV_X1 U79 ( .A(B[3]), .ZN(n101) );
  INV_X1 U80 ( .A(B[2]), .ZN(n102) );
  INV_X1 U81 ( .A(B[10]), .ZN(n94) );
  INV_X1 U82 ( .A(B[9]), .ZN(n95) );
  INV_X1 U83 ( .A(B[12]), .ZN(n92) );
  INV_X1 U84 ( .A(B[11]), .ZN(n93) );
  INV_X1 U85 ( .A(B[14]), .ZN(n90) );
  INV_X1 U86 ( .A(B[13]), .ZN(n91) );
  INV_X1 U87 ( .A(B[16]), .ZN(n88) );
  INV_X1 U88 ( .A(B[15]), .ZN(n89) );
  AND2_X1 U89 ( .A1(A[15]), .A2(SUMB_15__0_), .ZN(n68) );
  INV_X1 U90 ( .A(A[9]), .ZN(n77) );
  INV_X1 U91 ( .A(A[4]), .ZN(n82) );
  INV_X1 U92 ( .A(A[5]), .ZN(n81) );
  INV_X1 U93 ( .A(A[6]), .ZN(n80) );
  INV_X1 U94 ( .A(A[7]), .ZN(n79) );
  INV_X1 U95 ( .A(A[8]), .ZN(n78) );
  INV_X1 U96 ( .A(A[10]), .ZN(n76) );
  INV_X1 U97 ( .A(A[11]), .ZN(n75) );
  INV_X1 U98 ( .A(A[12]), .ZN(n74) );
  INV_X1 U99 ( .A(B[1]), .ZN(n103) );
  INV_X1 U100 ( .A(B[0]), .ZN(n104) );
  XOR2_X1 U101 ( .A(A[15]), .B(SUMB_15__0_), .Z(n69) );
  INV_X1 U102 ( .A(A[15]), .ZN(n71) );
  INV_X1 U103 ( .A(A[13]), .ZN(n73) );
  INV_X1 U104 ( .A(A[14]), .ZN(n72) );
  NOR2_X1 U105 ( .A1(n77), .A2(n95), .ZN(ab_9__9_) );
  NOR2_X1 U106 ( .A1(n77), .A2(n96), .ZN(ab_9__8_) );
  NOR2_X1 U107 ( .A1(n77), .A2(n97), .ZN(ab_9__7_) );
  NOR2_X1 U108 ( .A1(n77), .A2(n98), .ZN(ab_9__6_) );
  NOR2_X1 U109 ( .A1(n77), .A2(n99), .ZN(ab_9__5_) );
  NOR2_X1 U110 ( .A1(n77), .A2(n100), .ZN(ab_9__4_) );
  NOR2_X1 U111 ( .A1(n77), .A2(n101), .ZN(ab_9__3_) );
  NOR2_X1 U112 ( .A1(n77), .A2(n102), .ZN(ab_9__2_) );
  NOR2_X1 U113 ( .A1(n77), .A2(n103), .ZN(ab_9__1_) );
  NOR2_X1 U114 ( .A1(A[9]), .A2(n87), .ZN(ab_9__17_) );
  NOR2_X1 U115 ( .A1(n77), .A2(n88), .ZN(ab_9__16_) );
  NOR2_X1 U116 ( .A1(n77), .A2(n89), .ZN(ab_9__15_) );
  NOR2_X1 U117 ( .A1(n77), .A2(n90), .ZN(ab_9__14_) );
  NOR2_X1 U118 ( .A1(n77), .A2(n91), .ZN(ab_9__13_) );
  NOR2_X1 U119 ( .A1(n77), .A2(n92), .ZN(ab_9__12_) );
  NOR2_X1 U120 ( .A1(n77), .A2(n93), .ZN(ab_9__11_) );
  NOR2_X1 U121 ( .A1(n77), .A2(n94), .ZN(ab_9__10_) );
  NOR2_X1 U122 ( .A1(n77), .A2(n104), .ZN(ab_9__0_) );
  NOR2_X1 U123 ( .A1(n95), .A2(n78), .ZN(ab_8__9_) );
  NOR2_X1 U124 ( .A1(n96), .A2(n78), .ZN(ab_8__8_) );
  NOR2_X1 U125 ( .A1(n97), .A2(n78), .ZN(ab_8__7_) );
  NOR2_X1 U126 ( .A1(n98), .A2(n78), .ZN(ab_8__6_) );
  NOR2_X1 U127 ( .A1(n99), .A2(n78), .ZN(ab_8__5_) );
  NOR2_X1 U128 ( .A1(n100), .A2(n78), .ZN(ab_8__4_) );
  NOR2_X1 U129 ( .A1(n101), .A2(n78), .ZN(ab_8__3_) );
  NOR2_X1 U130 ( .A1(n102), .A2(n78), .ZN(ab_8__2_) );
  NOR2_X1 U131 ( .A1(n103), .A2(n78), .ZN(ab_8__1_) );
  NOR2_X1 U132 ( .A1(A[8]), .A2(n87), .ZN(ab_8__17_) );
  NOR2_X1 U133 ( .A1(n88), .A2(n78), .ZN(ab_8__16_) );
  NOR2_X1 U134 ( .A1(n89), .A2(n78), .ZN(ab_8__15_) );
  NOR2_X1 U135 ( .A1(n90), .A2(n78), .ZN(ab_8__14_) );
  NOR2_X1 U136 ( .A1(n91), .A2(n78), .ZN(ab_8__13_) );
  NOR2_X1 U137 ( .A1(n92), .A2(n78), .ZN(ab_8__12_) );
  NOR2_X1 U138 ( .A1(n93), .A2(n78), .ZN(ab_8__11_) );
  NOR2_X1 U139 ( .A1(n94), .A2(n78), .ZN(ab_8__10_) );
  NOR2_X1 U140 ( .A1(n104), .A2(n78), .ZN(ab_8__0_) );
  NOR2_X1 U141 ( .A1(n95), .A2(n79), .ZN(ab_7__9_) );
  NOR2_X1 U142 ( .A1(n96), .A2(n79), .ZN(ab_7__8_) );
  NOR2_X1 U143 ( .A1(n97), .A2(n79), .ZN(ab_7__7_) );
  NOR2_X1 U144 ( .A1(n98), .A2(n79), .ZN(ab_7__6_) );
  NOR2_X1 U145 ( .A1(n99), .A2(n79), .ZN(ab_7__5_) );
  NOR2_X1 U146 ( .A1(n100), .A2(n79), .ZN(ab_7__4_) );
  NOR2_X1 U147 ( .A1(n101), .A2(n79), .ZN(ab_7__3_) );
  NOR2_X1 U148 ( .A1(n102), .A2(n79), .ZN(ab_7__2_) );
  NOR2_X1 U149 ( .A1(n103), .A2(n79), .ZN(ab_7__1_) );
  NOR2_X1 U150 ( .A1(A[7]), .A2(n87), .ZN(ab_7__17_) );
  NOR2_X1 U151 ( .A1(n88), .A2(n79), .ZN(ab_7__16_) );
  NOR2_X1 U152 ( .A1(n89), .A2(n79), .ZN(ab_7__15_) );
  NOR2_X1 U153 ( .A1(n90), .A2(n79), .ZN(ab_7__14_) );
  NOR2_X1 U154 ( .A1(n91), .A2(n79), .ZN(ab_7__13_) );
  NOR2_X1 U155 ( .A1(n92), .A2(n79), .ZN(ab_7__12_) );
  NOR2_X1 U156 ( .A1(n93), .A2(n79), .ZN(ab_7__11_) );
  NOR2_X1 U157 ( .A1(n94), .A2(n79), .ZN(ab_7__10_) );
  NOR2_X1 U158 ( .A1(n104), .A2(n79), .ZN(ab_7__0_) );
  NOR2_X1 U159 ( .A1(n95), .A2(n80), .ZN(ab_6__9_) );
  NOR2_X1 U160 ( .A1(n96), .A2(n80), .ZN(ab_6__8_) );
  NOR2_X1 U161 ( .A1(n97), .A2(n80), .ZN(ab_6__7_) );
  NOR2_X1 U162 ( .A1(n98), .A2(n80), .ZN(ab_6__6_) );
  NOR2_X1 U163 ( .A1(n99), .A2(n80), .ZN(ab_6__5_) );
  NOR2_X1 U164 ( .A1(n100), .A2(n80), .ZN(ab_6__4_) );
  NOR2_X1 U165 ( .A1(n101), .A2(n80), .ZN(ab_6__3_) );
  NOR2_X1 U166 ( .A1(n102), .A2(n80), .ZN(ab_6__2_) );
  NOR2_X1 U167 ( .A1(n103), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U168 ( .A1(A[6]), .A2(n87), .ZN(ab_6__17_) );
  NOR2_X1 U169 ( .A1(n88), .A2(n80), .ZN(ab_6__16_) );
  NOR2_X1 U170 ( .A1(n89), .A2(n80), .ZN(ab_6__15_) );
  NOR2_X1 U171 ( .A1(n90), .A2(n80), .ZN(ab_6__14_) );
  NOR2_X1 U172 ( .A1(n91), .A2(n80), .ZN(ab_6__13_) );
  NOR2_X1 U173 ( .A1(n92), .A2(n80), .ZN(ab_6__12_) );
  NOR2_X1 U174 ( .A1(n93), .A2(n80), .ZN(ab_6__11_) );
  NOR2_X1 U175 ( .A1(n94), .A2(n80), .ZN(ab_6__10_) );
  NOR2_X1 U176 ( .A1(n104), .A2(n80), .ZN(ab_6__0_) );
  NOR2_X1 U177 ( .A1(n95), .A2(n81), .ZN(ab_5__9_) );
  NOR2_X1 U178 ( .A1(n96), .A2(n81), .ZN(ab_5__8_) );
  NOR2_X1 U179 ( .A1(n97), .A2(n81), .ZN(ab_5__7_) );
  NOR2_X1 U180 ( .A1(n98), .A2(n81), .ZN(ab_5__6_) );
  NOR2_X1 U181 ( .A1(n99), .A2(n81), .ZN(ab_5__5_) );
  NOR2_X1 U182 ( .A1(n100), .A2(n81), .ZN(ab_5__4_) );
  NOR2_X1 U183 ( .A1(n101), .A2(n81), .ZN(ab_5__3_) );
  NOR2_X1 U184 ( .A1(n102), .A2(n81), .ZN(ab_5__2_) );
  NOR2_X1 U185 ( .A1(n103), .A2(n81), .ZN(ab_5__1_) );
  NOR2_X1 U186 ( .A1(A[5]), .A2(n87), .ZN(ab_5__17_) );
  NOR2_X1 U187 ( .A1(n88), .A2(n81), .ZN(ab_5__16_) );
  NOR2_X1 U188 ( .A1(n89), .A2(n81), .ZN(ab_5__15_) );
  NOR2_X1 U189 ( .A1(n90), .A2(n81), .ZN(ab_5__14_) );
  NOR2_X1 U190 ( .A1(n91), .A2(n81), .ZN(ab_5__13_) );
  NOR2_X1 U191 ( .A1(n92), .A2(n81), .ZN(ab_5__12_) );
  NOR2_X1 U192 ( .A1(n93), .A2(n81), .ZN(ab_5__11_) );
  NOR2_X1 U193 ( .A1(n94), .A2(n81), .ZN(ab_5__10_) );
  NOR2_X1 U194 ( .A1(n104), .A2(n81), .ZN(ab_5__0_) );
  NOR2_X1 U195 ( .A1(n95), .A2(n82), .ZN(ab_4__9_) );
  NOR2_X1 U196 ( .A1(n96), .A2(n82), .ZN(ab_4__8_) );
  NOR2_X1 U197 ( .A1(n97), .A2(n82), .ZN(ab_4__7_) );
  NOR2_X1 U198 ( .A1(n98), .A2(n82), .ZN(ab_4__6_) );
  NOR2_X1 U199 ( .A1(n99), .A2(n82), .ZN(ab_4__5_) );
  NOR2_X1 U200 ( .A1(n100), .A2(n82), .ZN(ab_4__4_) );
  NOR2_X1 U201 ( .A1(n101), .A2(n82), .ZN(ab_4__3_) );
  NOR2_X1 U202 ( .A1(n102), .A2(n82), .ZN(ab_4__2_) );
  NOR2_X1 U203 ( .A1(n103), .A2(n82), .ZN(ab_4__1_) );
  NOR2_X1 U204 ( .A1(A[4]), .A2(n87), .ZN(ab_4__17_) );
  NOR2_X1 U205 ( .A1(n88), .A2(n82), .ZN(ab_4__16_) );
  NOR2_X1 U206 ( .A1(n89), .A2(n82), .ZN(ab_4__15_) );
  NOR2_X1 U207 ( .A1(n90), .A2(n82), .ZN(ab_4__14_) );
  NOR2_X1 U208 ( .A1(n91), .A2(n82), .ZN(ab_4__13_) );
  NOR2_X1 U209 ( .A1(n92), .A2(n82), .ZN(ab_4__12_) );
  NOR2_X1 U210 ( .A1(n93), .A2(n82), .ZN(ab_4__11_) );
  NOR2_X1 U211 ( .A1(n94), .A2(n82), .ZN(ab_4__10_) );
  NOR2_X1 U212 ( .A1(n104), .A2(n82), .ZN(ab_4__0_) );
  NOR2_X1 U213 ( .A1(n95), .A2(n83), .ZN(ab_3__9_) );
  NOR2_X1 U214 ( .A1(n96), .A2(n83), .ZN(ab_3__8_) );
  NOR2_X1 U215 ( .A1(n97), .A2(n83), .ZN(ab_3__7_) );
  NOR2_X1 U216 ( .A1(n98), .A2(n83), .ZN(ab_3__6_) );
  NOR2_X1 U217 ( .A1(n99), .A2(n83), .ZN(ab_3__5_) );
  NOR2_X1 U218 ( .A1(n100), .A2(n83), .ZN(ab_3__4_) );
  NOR2_X1 U219 ( .A1(n101), .A2(n83), .ZN(ab_3__3_) );
  NOR2_X1 U220 ( .A1(n102), .A2(n83), .ZN(ab_3__2_) );
  NOR2_X1 U221 ( .A1(n103), .A2(n83), .ZN(ab_3__1_) );
  NOR2_X1 U222 ( .A1(A[3]), .A2(n87), .ZN(ab_3__17_) );
  NOR2_X1 U223 ( .A1(n88), .A2(n83), .ZN(ab_3__16_) );
  NOR2_X1 U224 ( .A1(n89), .A2(n83), .ZN(ab_3__15_) );
  NOR2_X1 U225 ( .A1(n90), .A2(n83), .ZN(ab_3__14_) );
  NOR2_X1 U226 ( .A1(n91), .A2(n83), .ZN(ab_3__13_) );
  NOR2_X1 U227 ( .A1(n92), .A2(n83), .ZN(ab_3__12_) );
  NOR2_X1 U228 ( .A1(n93), .A2(n83), .ZN(ab_3__11_) );
  NOR2_X1 U229 ( .A1(n94), .A2(n83), .ZN(ab_3__10_) );
  NOR2_X1 U230 ( .A1(n104), .A2(n83), .ZN(ab_3__0_) );
  NOR2_X1 U231 ( .A1(n95), .A2(n84), .ZN(ab_2__9_) );
  NOR2_X1 U232 ( .A1(n96), .A2(n84), .ZN(ab_2__8_) );
  NOR2_X1 U233 ( .A1(n97), .A2(n84), .ZN(ab_2__7_) );
  NOR2_X1 U234 ( .A1(n98), .A2(n84), .ZN(ab_2__6_) );
  NOR2_X1 U235 ( .A1(n99), .A2(n84), .ZN(ab_2__5_) );
  NOR2_X1 U236 ( .A1(n100), .A2(n84), .ZN(ab_2__4_) );
  NOR2_X1 U237 ( .A1(n101), .A2(n84), .ZN(ab_2__3_) );
  NOR2_X1 U238 ( .A1(n102), .A2(n84), .ZN(ab_2__2_) );
  NOR2_X1 U239 ( .A1(n103), .A2(n84), .ZN(ab_2__1_) );
  NOR2_X1 U240 ( .A1(A[2]), .A2(n87), .ZN(ab_2__17_) );
  NOR2_X1 U241 ( .A1(n88), .A2(n84), .ZN(ab_2__16_) );
  NOR2_X1 U242 ( .A1(n89), .A2(n84), .ZN(ab_2__15_) );
  NOR2_X1 U243 ( .A1(n90), .A2(n84), .ZN(ab_2__14_) );
  NOR2_X1 U244 ( .A1(n91), .A2(n84), .ZN(ab_2__13_) );
  NOR2_X1 U245 ( .A1(n92), .A2(n84), .ZN(ab_2__12_) );
  NOR2_X1 U246 ( .A1(n93), .A2(n84), .ZN(ab_2__11_) );
  NOR2_X1 U247 ( .A1(n94), .A2(n84), .ZN(ab_2__10_) );
  NOR2_X1 U248 ( .A1(n104), .A2(n84), .ZN(ab_2__0_) );
  NOR2_X1 U249 ( .A1(n95), .A2(n85), .ZN(ab_1__9_) );
  NOR2_X1 U250 ( .A1(n96), .A2(n85), .ZN(ab_1__8_) );
  NOR2_X1 U251 ( .A1(n97), .A2(n85), .ZN(ab_1__7_) );
  NOR2_X1 U252 ( .A1(n98), .A2(n85), .ZN(ab_1__6_) );
  NOR2_X1 U253 ( .A1(n99), .A2(n85), .ZN(ab_1__5_) );
  NOR2_X1 U254 ( .A1(n100), .A2(n85), .ZN(ab_1__4_) );
  NOR2_X1 U255 ( .A1(n101), .A2(n85), .ZN(ab_1__3_) );
  NOR2_X1 U256 ( .A1(n102), .A2(n85), .ZN(ab_1__2_) );
  NOR2_X1 U257 ( .A1(n103), .A2(n85), .ZN(ab_1__1_) );
  NOR2_X1 U258 ( .A1(A[1]), .A2(n87), .ZN(ab_1__17_) );
  NOR2_X1 U259 ( .A1(n88), .A2(n85), .ZN(ab_1__16_) );
  NOR2_X1 U260 ( .A1(n89), .A2(n85), .ZN(ab_1__15_) );
  NOR2_X1 U261 ( .A1(n90), .A2(n85), .ZN(ab_1__14_) );
  NOR2_X1 U262 ( .A1(n91), .A2(n85), .ZN(ab_1__13_) );
  NOR2_X1 U263 ( .A1(n92), .A2(n85), .ZN(ab_1__12_) );
  NOR2_X1 U264 ( .A1(n93), .A2(n85), .ZN(ab_1__11_) );
  NOR2_X1 U265 ( .A1(n94), .A2(n85), .ZN(ab_1__10_) );
  NOR2_X1 U266 ( .A1(n104), .A2(n85), .ZN(ab_1__0_) );
  NOR2_X1 U267 ( .A1(B[9]), .A2(n71), .ZN(ab_15__9_) );
  NOR2_X1 U268 ( .A1(B[8]), .A2(n71), .ZN(ab_15__8_) );
  NOR2_X1 U269 ( .A1(B[7]), .A2(n71), .ZN(ab_15__7_) );
  NOR2_X1 U270 ( .A1(B[6]), .A2(n71), .ZN(ab_15__6_) );
  NOR2_X1 U271 ( .A1(B[5]), .A2(n71), .ZN(ab_15__5_) );
  NOR2_X1 U272 ( .A1(B[4]), .A2(n71), .ZN(ab_15__4_) );
  NOR2_X1 U273 ( .A1(B[3]), .A2(n71), .ZN(ab_15__3_) );
  NOR2_X1 U274 ( .A1(B[2]), .A2(n71), .ZN(ab_15__2_) );
  NOR2_X1 U275 ( .A1(B[1]), .A2(n71), .ZN(ab_15__1_) );
  NOR2_X1 U276 ( .A1(n87), .A2(n71), .ZN(ab_15__17_) );
  NOR2_X1 U277 ( .A1(B[16]), .A2(n71), .ZN(ab_15__16_) );
  NOR2_X1 U278 ( .A1(B[15]), .A2(n71), .ZN(ab_15__15_) );
  NOR2_X1 U279 ( .A1(B[14]), .A2(n71), .ZN(ab_15__14_) );
  NOR2_X1 U280 ( .A1(B[13]), .A2(n71), .ZN(ab_15__13_) );
  NOR2_X1 U281 ( .A1(B[12]), .A2(n71), .ZN(ab_15__12_) );
  NOR2_X1 U282 ( .A1(B[11]), .A2(n71), .ZN(ab_15__11_) );
  NOR2_X1 U283 ( .A1(B[10]), .A2(n71), .ZN(ab_15__10_) );
  NOR2_X1 U284 ( .A1(B[0]), .A2(n71), .ZN(ab_15__0_) );
  NOR2_X1 U285 ( .A1(n95), .A2(n72), .ZN(ab_14__9_) );
  NOR2_X1 U286 ( .A1(n96), .A2(n72), .ZN(ab_14__8_) );
  NOR2_X1 U287 ( .A1(n97), .A2(n72), .ZN(ab_14__7_) );
  NOR2_X1 U288 ( .A1(n98), .A2(n72), .ZN(ab_14__6_) );
  NOR2_X1 U289 ( .A1(n99), .A2(n72), .ZN(ab_14__5_) );
  NOR2_X1 U290 ( .A1(n100), .A2(n72), .ZN(ab_14__4_) );
  NOR2_X1 U291 ( .A1(n101), .A2(n72), .ZN(ab_14__3_) );
  NOR2_X1 U292 ( .A1(n102), .A2(n72), .ZN(ab_14__2_) );
  NOR2_X1 U293 ( .A1(n103), .A2(n72), .ZN(ab_14__1_) );
  NOR2_X1 U294 ( .A1(A[14]), .A2(n87), .ZN(ab_14__17_) );
  NOR2_X1 U295 ( .A1(n88), .A2(n72), .ZN(ab_14__16_) );
  NOR2_X1 U296 ( .A1(n89), .A2(n72), .ZN(ab_14__15_) );
  NOR2_X1 U297 ( .A1(n90), .A2(n72), .ZN(ab_14__14_) );
  NOR2_X1 U298 ( .A1(n91), .A2(n72), .ZN(ab_14__13_) );
  NOR2_X1 U299 ( .A1(n92), .A2(n72), .ZN(ab_14__12_) );
  NOR2_X1 U300 ( .A1(n93), .A2(n72), .ZN(ab_14__11_) );
  NOR2_X1 U301 ( .A1(n94), .A2(n72), .ZN(ab_14__10_) );
  NOR2_X1 U302 ( .A1(n104), .A2(n72), .ZN(ab_14__0_) );
  NOR2_X1 U303 ( .A1(n95), .A2(n73), .ZN(ab_13__9_) );
  NOR2_X1 U304 ( .A1(n96), .A2(n73), .ZN(ab_13__8_) );
  NOR2_X1 U305 ( .A1(n97), .A2(n73), .ZN(ab_13__7_) );
  NOR2_X1 U306 ( .A1(n98), .A2(n73), .ZN(ab_13__6_) );
  NOR2_X1 U307 ( .A1(n99), .A2(n73), .ZN(ab_13__5_) );
  NOR2_X1 U308 ( .A1(n100), .A2(n73), .ZN(ab_13__4_) );
  NOR2_X1 U309 ( .A1(n101), .A2(n73), .ZN(ab_13__3_) );
  NOR2_X1 U310 ( .A1(n102), .A2(n73), .ZN(ab_13__2_) );
  NOR2_X1 U311 ( .A1(n103), .A2(n73), .ZN(ab_13__1_) );
  NOR2_X1 U312 ( .A1(A[13]), .A2(n87), .ZN(ab_13__17_) );
  NOR2_X1 U313 ( .A1(n88), .A2(n73), .ZN(ab_13__16_) );
  NOR2_X1 U314 ( .A1(n89), .A2(n73), .ZN(ab_13__15_) );
  NOR2_X1 U315 ( .A1(n90), .A2(n73), .ZN(ab_13__14_) );
  NOR2_X1 U316 ( .A1(n91), .A2(n73), .ZN(ab_13__13_) );
  NOR2_X1 U317 ( .A1(n92), .A2(n73), .ZN(ab_13__12_) );
  NOR2_X1 U318 ( .A1(n93), .A2(n73), .ZN(ab_13__11_) );
  NOR2_X1 U319 ( .A1(n94), .A2(n73), .ZN(ab_13__10_) );
  NOR2_X1 U320 ( .A1(n104), .A2(n73), .ZN(ab_13__0_) );
  NOR2_X1 U321 ( .A1(n95), .A2(n74), .ZN(ab_12__9_) );
  NOR2_X1 U322 ( .A1(n96), .A2(n74), .ZN(ab_12__8_) );
  NOR2_X1 U323 ( .A1(n97), .A2(n74), .ZN(ab_12__7_) );
  NOR2_X1 U324 ( .A1(n98), .A2(n74), .ZN(ab_12__6_) );
  NOR2_X1 U325 ( .A1(n99), .A2(n74), .ZN(ab_12__5_) );
  NOR2_X1 U326 ( .A1(n100), .A2(n74), .ZN(ab_12__4_) );
  NOR2_X1 U327 ( .A1(n101), .A2(n74), .ZN(ab_12__3_) );
  NOR2_X1 U328 ( .A1(n102), .A2(n74), .ZN(ab_12__2_) );
  NOR2_X1 U329 ( .A1(n103), .A2(n74), .ZN(ab_12__1_) );
  NOR2_X1 U330 ( .A1(A[12]), .A2(n87), .ZN(ab_12__17_) );
  NOR2_X1 U331 ( .A1(n88), .A2(n74), .ZN(ab_12__16_) );
  NOR2_X1 U332 ( .A1(n89), .A2(n74), .ZN(ab_12__15_) );
  NOR2_X1 U333 ( .A1(n90), .A2(n74), .ZN(ab_12__14_) );
  NOR2_X1 U334 ( .A1(n91), .A2(n74), .ZN(ab_12__13_) );
  NOR2_X1 U335 ( .A1(n92), .A2(n74), .ZN(ab_12__12_) );
  NOR2_X1 U336 ( .A1(n93), .A2(n74), .ZN(ab_12__11_) );
  NOR2_X1 U337 ( .A1(n94), .A2(n74), .ZN(ab_12__10_) );
  NOR2_X1 U338 ( .A1(n104), .A2(n74), .ZN(ab_12__0_) );
  NOR2_X1 U339 ( .A1(n95), .A2(n75), .ZN(ab_11__9_) );
  NOR2_X1 U340 ( .A1(n96), .A2(n75), .ZN(ab_11__8_) );
  NOR2_X1 U341 ( .A1(n97), .A2(n75), .ZN(ab_11__7_) );
  NOR2_X1 U342 ( .A1(n98), .A2(n75), .ZN(ab_11__6_) );
  NOR2_X1 U343 ( .A1(n99), .A2(n75), .ZN(ab_11__5_) );
  NOR2_X1 U344 ( .A1(n100), .A2(n75), .ZN(ab_11__4_) );
  NOR2_X1 U345 ( .A1(n101), .A2(n75), .ZN(ab_11__3_) );
  NOR2_X1 U346 ( .A1(n102), .A2(n75), .ZN(ab_11__2_) );
  NOR2_X1 U347 ( .A1(n103), .A2(n75), .ZN(ab_11__1_) );
  NOR2_X1 U348 ( .A1(A[11]), .A2(n87), .ZN(ab_11__17_) );
  NOR2_X1 U349 ( .A1(n88), .A2(n75), .ZN(ab_11__16_) );
  NOR2_X1 U350 ( .A1(n89), .A2(n75), .ZN(ab_11__15_) );
  NOR2_X1 U351 ( .A1(n90), .A2(n75), .ZN(ab_11__14_) );
  NOR2_X1 U352 ( .A1(n91), .A2(n75), .ZN(ab_11__13_) );
  NOR2_X1 U353 ( .A1(n92), .A2(n75), .ZN(ab_11__12_) );
  NOR2_X1 U354 ( .A1(n93), .A2(n75), .ZN(ab_11__11_) );
  NOR2_X1 U355 ( .A1(n94), .A2(n75), .ZN(ab_11__10_) );
  NOR2_X1 U356 ( .A1(n104), .A2(n75), .ZN(ab_11__0_) );
  NOR2_X1 U357 ( .A1(n95), .A2(n76), .ZN(ab_10__9_) );
  NOR2_X1 U358 ( .A1(n96), .A2(n76), .ZN(ab_10__8_) );
  NOR2_X1 U359 ( .A1(n97), .A2(n76), .ZN(ab_10__7_) );
  NOR2_X1 U360 ( .A1(n98), .A2(n76), .ZN(ab_10__6_) );
  NOR2_X1 U361 ( .A1(n99), .A2(n76), .ZN(ab_10__5_) );
  NOR2_X1 U362 ( .A1(n100), .A2(n76), .ZN(ab_10__4_) );
  NOR2_X1 U363 ( .A1(n101), .A2(n76), .ZN(ab_10__3_) );
  NOR2_X1 U364 ( .A1(n102), .A2(n76), .ZN(ab_10__2_) );
  NOR2_X1 U365 ( .A1(n103), .A2(n76), .ZN(ab_10__1_) );
  NOR2_X1 U366 ( .A1(A[10]), .A2(n87), .ZN(ab_10__17_) );
  NOR2_X1 U367 ( .A1(n88), .A2(n76), .ZN(ab_10__16_) );
  NOR2_X1 U368 ( .A1(n89), .A2(n76), .ZN(ab_10__15_) );
  NOR2_X1 U369 ( .A1(n90), .A2(n76), .ZN(ab_10__14_) );
  NOR2_X1 U370 ( .A1(n91), .A2(n76), .ZN(ab_10__13_) );
  NOR2_X1 U371 ( .A1(n92), .A2(n76), .ZN(ab_10__12_) );
  NOR2_X1 U372 ( .A1(n93), .A2(n76), .ZN(ab_10__11_) );
  NOR2_X1 U373 ( .A1(n94), .A2(n76), .ZN(ab_10__10_) );
  NOR2_X1 U374 ( .A1(n104), .A2(n76), .ZN(ab_10__0_) );
  NOR2_X1 U375 ( .A1(n95), .A2(n86), .ZN(ab_0__9_) );
  NOR2_X1 U376 ( .A1(n96), .A2(n86), .ZN(ab_0__8_) );
  NOR2_X1 U377 ( .A1(n97), .A2(n86), .ZN(ab_0__7_) );
  NOR2_X1 U378 ( .A1(n98), .A2(n86), .ZN(ab_0__6_) );
  NOR2_X1 U379 ( .A1(n99), .A2(n86), .ZN(ab_0__5_) );
  NOR2_X1 U380 ( .A1(n100), .A2(n86), .ZN(ab_0__4_) );
  NOR2_X1 U381 ( .A1(n101), .A2(n86), .ZN(ab_0__3_) );
  NOR2_X1 U382 ( .A1(n102), .A2(n86), .ZN(ab_0__2_) );
  NOR2_X1 U383 ( .A1(n103), .A2(n86), .ZN(ab_0__1_) );
  NOR2_X1 U384 ( .A1(A[0]), .A2(n87), .ZN(ab_0__17_) );
  NOR2_X1 U385 ( .A1(n88), .A2(n86), .ZN(ab_0__16_) );
  NOR2_X1 U386 ( .A1(n89), .A2(n86), .ZN(ab_0__15_) );
  NOR2_X1 U387 ( .A1(n90), .A2(n86), .ZN(ab_0__14_) );
  NOR2_X1 U388 ( .A1(n91), .A2(n86), .ZN(ab_0__13_) );
  NOR2_X1 U389 ( .A1(n92), .A2(n86), .ZN(ab_0__12_) );
  NOR2_X1 U390 ( .A1(n93), .A2(n86), .ZN(ab_0__11_) );
  NOR2_X1 U391 ( .A1(n94), .A2(n86), .ZN(ab_0__10_) );
  NOR2_X1 U392 ( .A1(n104), .A2(n86), .ZN(PRODUCT[0]) );
endmodule


module gng_smul_16_18 ( clk, a, b, p );
  input [15:0] a;
  input [17:0] b;
  output [33:0] p;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33;
  wire   [15:0] a_reg;
  wire   [17:0] b_reg;

  DFF_X1 a_reg_reg_15_ ( .D(a[15]), .CK(clk), .Q(a_reg[15]) );
  DFF_X1 a_reg_reg_14_ ( .D(a[14]), .CK(clk), .Q(a_reg[14]) );
  DFF_X1 a_reg_reg_13_ ( .D(a[13]), .CK(clk), .Q(a_reg[13]) );
  DFF_X1 a_reg_reg_12_ ( .D(a[12]), .CK(clk), .Q(a_reg[12]) );
  DFF_X1 a_reg_reg_11_ ( .D(a[11]), .CK(clk), .Q(a_reg[11]) );
  DFF_X1 a_reg_reg_10_ ( .D(a[10]), .CK(clk), .Q(a_reg[10]) );
  DFF_X1 a_reg_reg_9_ ( .D(a[9]), .CK(clk), .Q(a_reg[9]) );
  DFF_X1 a_reg_reg_8_ ( .D(a[8]), .CK(clk), .Q(a_reg[8]) );
  DFF_X1 a_reg_reg_7_ ( .D(a[7]), .CK(clk), .Q(a_reg[7]) );
  DFF_X1 a_reg_reg_6_ ( .D(a[6]), .CK(clk), .Q(a_reg[6]) );
  DFF_X1 a_reg_reg_5_ ( .D(a[5]), .CK(clk), .Q(a_reg[5]) );
  DFF_X1 a_reg_reg_4_ ( .D(a[4]), .CK(clk), .Q(a_reg[4]) );
  DFF_X1 a_reg_reg_3_ ( .D(a[3]), .CK(clk), .Q(a_reg[3]) );
  DFF_X1 a_reg_reg_2_ ( .D(a[2]), .CK(clk), .Q(a_reg[2]) );
  DFF_X1 a_reg_reg_1_ ( .D(a[1]), .CK(clk), .Q(a_reg[1]) );
  DFF_X1 a_reg_reg_0_ ( .D(a[0]), .CK(clk), .Q(a_reg[0]) );
  DFF_X1 b_reg_reg_17_ ( .D(b[17]), .CK(clk), .Q(b_reg[17]) );
  DFF_X1 b_reg_reg_16_ ( .D(b[16]), .CK(clk), .Q(b_reg[16]) );
  DFF_X1 b_reg_reg_15_ ( .D(b[15]), .CK(clk), .Q(b_reg[15]) );
  DFF_X1 b_reg_reg_14_ ( .D(b[14]), .CK(clk), .Q(b_reg[14]) );
  DFF_X1 b_reg_reg_13_ ( .D(b[13]), .CK(clk), .Q(b_reg[13]) );
  DFF_X1 b_reg_reg_12_ ( .D(b[12]), .CK(clk), .Q(b_reg[12]) );
  DFF_X1 b_reg_reg_11_ ( .D(b[11]), .CK(clk), .Q(b_reg[11]) );
  DFF_X1 b_reg_reg_10_ ( .D(b[10]), .CK(clk), .Q(b_reg[10]) );
  DFF_X1 b_reg_reg_9_ ( .D(b[9]), .CK(clk), .Q(b_reg[9]) );
  DFF_X1 b_reg_reg_8_ ( .D(b[8]), .CK(clk), .Q(b_reg[8]) );
  DFF_X1 b_reg_reg_7_ ( .D(b[7]), .CK(clk), .Q(b_reg[7]) );
  DFF_X1 b_reg_reg_6_ ( .D(b[6]), .CK(clk), .Q(b_reg[6]) );
  DFF_X1 b_reg_reg_5_ ( .D(b[5]), .CK(clk), .Q(b_reg[5]) );
  DFF_X1 b_reg_reg_4_ ( .D(b[4]), .CK(clk), .Q(b_reg[4]) );
  DFF_X1 b_reg_reg_3_ ( .D(b[3]), .CK(clk), .Q(b_reg[3]) );
  DFF_X1 b_reg_reg_2_ ( .D(b[2]), .CK(clk), .Q(b_reg[2]) );
  DFF_X1 b_reg_reg_1_ ( .D(b[1]), .CK(clk), .Q(b_reg[1]) );
  DFF_X1 b_reg_reg_0_ ( .D(b[0]), .CK(clk), .Q(b_reg[0]) );
  DFF_X1 prod_reg_33_ ( .D(N33), .CK(clk), .Q(p[33]) );
  DFF_X1 prod_reg_32_ ( .D(N32), .CK(clk), .Q(p[32]) );
  DFF_X1 prod_reg_31_ ( .D(N31), .CK(clk), .Q(p[31]) );
  DFF_X1 prod_reg_30_ ( .D(N30), .CK(clk), .Q(p[30]) );
  DFF_X1 prod_reg_29_ ( .D(N29), .CK(clk), .Q(p[29]) );
  DFF_X1 prod_reg_28_ ( .D(N28), .CK(clk), .Q(p[28]) );
  DFF_X1 prod_reg_27_ ( .D(N27), .CK(clk), .Q(p[27]) );
  DFF_X1 prod_reg_26_ ( .D(N26), .CK(clk), .Q(p[26]) );
  DFF_X1 prod_reg_25_ ( .D(N25), .CK(clk), .Q(p[25]) );
  DFF_X1 prod_reg_24_ ( .D(N24), .CK(clk), .Q(p[24]) );
  DFF_X1 prod_reg_23_ ( .D(N23), .CK(clk), .Q(p[23]) );
  DFF_X1 prod_reg_22_ ( .D(N22), .CK(clk), .Q(p[22]) );
  DFF_X1 prod_reg_21_ ( .D(N21), .CK(clk), .Q(p[21]) );
  DFF_X1 prod_reg_20_ ( .D(N20), .CK(clk), .Q(p[20]) );
  DFF_X1 prod_reg_19_ ( .D(N19), .CK(clk), .Q(p[19]) );
  DFF_X1 prod_reg_18_ ( .D(N18), .CK(clk), .Q(p[18]) );
  DFF_X1 prod_reg_17_ ( .D(N17), .CK(clk), .Q(p[17]) );
  DFF_X1 prod_reg_16_ ( .D(N16), .CK(clk), .Q(p[16]) );
  DFF_X1 prod_reg_15_ ( .D(N15), .CK(clk), .Q(p[15]) );
  DFF_X1 prod_reg_14_ ( .D(N14), .CK(clk), .Q(p[14]) );
  DFF_X1 prod_reg_13_ ( .D(N13), .CK(clk), .Q(p[13]) );
  DFF_X1 prod_reg_12_ ( .D(N12), .CK(clk), .Q(p[12]) );
  DFF_X1 prod_reg_11_ ( .D(N11), .CK(clk), .Q(p[11]) );
  DFF_X1 prod_reg_10_ ( .D(N10), .CK(clk), .Q(p[10]) );
  DFF_X1 prod_reg_9_ ( .D(N9), .CK(clk), .Q(p[9]) );
  DFF_X1 prod_reg_8_ ( .D(N8), .CK(clk), .Q(p[8]) );
  DFF_X1 prod_reg_7_ ( .D(N7), .CK(clk), .Q(p[7]) );
  DFF_X1 prod_reg_6_ ( .D(N6), .CK(clk), .Q(p[6]) );
  DFF_X1 prod_reg_5_ ( .D(N5), .CK(clk), .Q(p[5]) );
  DFF_X1 prod_reg_4_ ( .D(N4), .CK(clk), .Q(p[4]) );
  DFF_X1 prod_reg_3_ ( .D(N3), .CK(clk), .Q(p[3]) );
  DFF_X1 prod_reg_2_ ( .D(N2), .CK(clk), .Q(p[2]) );
  DFF_X1 prod_reg_1_ ( .D(N1), .CK(clk), .Q(p[1]) );
  DFF_X1 prod_reg_0_ ( .D(N0), .CK(clk), .Q(p[0]) );
  gng_smul_16_18_DW02_mult_0 mult_60 ( .A(a_reg), .B(b_reg), .TC(1'b1), 
        .PRODUCT({N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4, N3, N2, N1, N0}) );
endmodule


module gng_interp_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(carry[15]), .ZN(SUM[15]) );
endmodule


module gng_interp_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [17:2] carry;

  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .S(SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INV_X1 U1 ( .A(A[1]), .ZN(n2) );
  INV_X1 U2 ( .A(B[1]), .ZN(n1) );
  OAI21_X1 U3 ( .B1(n2), .B2(n1), .A(n3), .ZN(carry[2]) );
  OAI211_X1 U4 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n3) );
endmodule


module gng_interp ( clk, rstn, valid_in, data_in, valid_out, data_out );
  input [63:0] data_in;
  output [15:0] data_out;
  input clk, rstn, valid_in;
  output valid_out;
  wire   N6, N7, N8, N9, N10, N11, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, N147, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         n710, n810, n910, n1010, n1110, n12, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n1, n3, n4, n5, n610, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n57, n58, n59, n600, n611, n620, n630, n640, n650, n660, n670,
         n680, n690, n700, n711, n720, n730, n740, n750, n760, n770, n780,
         n790, n800, n811, n820, n830, n840, n850, n860, n870, n880, n890,
         n900, n911, n920, n930, n940, n950, n960, n970, n980, n990, n1000,
         n1011, n1020, n1030, n1040, n1050, n1060, n1070, n1080, n1090, n1100,
         n1111, n1120, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43;
  wire   [5:0] num_lzd;
  wire   [5:0] num_lzd_r;
  wire   [1:0] offset;
  wire   [17:0] c0;
  wire   [17:0] c1;
  wire   [16:0] c2;
  wire   [14:0] x_r1;
  wire   [14:0] x_r2;
  wire   [14:0] x_r4;
  wire   [14:0] x_r3;
  wire   [17:0] c1_r1;
  wire   [17:0] c0_r1;
  wire   [17:0] c0_r2;
  wire   [17:0] c0_r3;
  wire   [17:0] c0_r5;
  wire   [17:0] c0_r4;
  wire   [8:0] sign_r;
  wire   [8:0] valid_in_r;
  wire   [37:20] sum1;
  wire   [32:19] mul1;
  wire   [16:2] sum2;

  DFF_X1 num_lzd_r_reg_5_ ( .D(N11), .CK(clk), .Q(num_lzd_r[5]) );
  DFF_X1 num_lzd_r_reg_4_ ( .D(N10), .CK(clk), .Q(num_lzd_r[4]), .QN(n710) );
  DFF_X1 num_lzd_r_reg_3_ ( .D(N9), .CK(clk), .Q(num_lzd_r[3]), .QN(n810) );
  DFF_X1 num_lzd_r_reg_2_ ( .D(N8), .CK(clk), .Q(num_lzd_r[2]), .QN(n910) );
  DFF_X1 num_lzd_r_reg_1_ ( .D(N7), .CK(clk), .Q(num_lzd_r[1]), .QN(n1010) );
  DFF_X1 num_lzd_r_reg_0_ ( .D(N6), .CK(clk), .Q(num_lzd_r[0]), .QN(n1110) );
  DFF_X1 mask_reg_14_ ( .D(N74), .CK(clk), .QN(n880) );
  DFF_X1 mask_reg_13_ ( .D(N73), .CK(clk), .QN(n860) );
  DFF_X1 mask_reg_12_ ( .D(N72), .CK(clk), .QN(n840) );
  DFF_X1 mask_reg_11_ ( .D(N71), .CK(clk), .QN(n820) );
  DFF_X1 mask_reg_10_ ( .D(N70), .CK(clk), .QN(n800) );
  DFF_X1 mask_reg_9_ ( .D(N69), .CK(clk), .QN(n780) );
  DFF_X1 mask_reg_8_ ( .D(N68), .CK(clk), .QN(n760) );
  DFF_X1 mask_reg_7_ ( .D(N67), .CK(clk), .QN(n740) );
  DFF_X1 mask_reg_6_ ( .D(N66), .CK(clk), .QN(n720) );
  DFF_X1 mask_reg_5_ ( .D(N65), .CK(clk), .QN(n700) );
  DFF_X1 mask_reg_4_ ( .D(N64), .CK(clk), .QN(n680) );
  DFF_X1 mask_reg_3_ ( .D(N63), .CK(clk), .QN(n660) );
  DFF_X1 mask_reg_2_ ( .D(N62), .CK(clk), .QN(n640) );
  DFF_X1 mask_reg_1_ ( .D(N61), .CK(clk), .QN(n620) );
  DFF_X1 mask_reg_0_ ( .D(N60), .CK(clk), .QN(n600) );
  DFF_X1 offset_reg_1_ ( .D(N76), .CK(clk), .Q(offset[1]) );
  DFF_X1 offset_reg_0_ ( .D(N75), .CK(clk), .Q(offset[0]) );
  DFF_X1 x_reg_14_ ( .D(N91), .CK(clk), .QN(n870) );
  DFF_X1 x_reg_13_ ( .D(N90), .CK(clk), .QN(n850) );
  DFF_X1 x_reg_12_ ( .D(N89), .CK(clk), .QN(n830) );
  DFF_X1 x_reg_11_ ( .D(N88), .CK(clk), .QN(n811) );
  DFF_X1 x_reg_10_ ( .D(N87), .CK(clk), .QN(n790) );
  DFF_X1 x_reg_9_ ( .D(N86), .CK(clk), .QN(n770) );
  DFF_X1 x_reg_8_ ( .D(N85), .CK(clk), .QN(n750) );
  DFF_X1 x_reg_7_ ( .D(N84), .CK(clk), .QN(n730) );
  DFF_X1 x_reg_6_ ( .D(N83), .CK(clk), .QN(n711) );
  DFF_X1 x_reg_5_ ( .D(N82), .CK(clk), .QN(n690) );
  DFF_X1 x_reg_4_ ( .D(N81), .CK(clk), .QN(n670) );
  DFF_X1 x_reg_3_ ( .D(N80), .CK(clk), .QN(n650) );
  DFF_X1 x_reg_2_ ( .D(N79), .CK(clk), .QN(n630) );
  DFF_X1 x_reg_1_ ( .D(N78), .CK(clk), .QN(n611) );
  DFF_X1 x_reg_0_ ( .D(N77), .CK(clk), .QN(n59) );
  DFF_X1 x_r1_reg_14_ ( .D(N92), .CK(clk), .Q(x_r1[14]) );
  DFF_X1 x_r2_reg_14_ ( .D(x_r1[14]), .CK(clk), .Q(x_r2[14]) );
  DFF_X1 x_r3_reg_14_ ( .D(x_r2[14]), .CK(clk), .Q(x_r3[14]) );
  DFF_X1 x_r1_reg_13_ ( .D(N93), .CK(clk), .Q(x_r1[13]) );
  DFF_X1 x_r2_reg_13_ ( .D(x_r1[13]), .CK(clk), .Q(x_r2[13]) );
  DFF_X1 x_r3_reg_13_ ( .D(x_r2[13]), .CK(clk), .Q(x_r3[13]) );
  DFF_X1 x_r1_reg_12_ ( .D(N94), .CK(clk), .Q(x_r1[12]) );
  DFF_X1 x_r2_reg_12_ ( .D(x_r1[12]), .CK(clk), .Q(x_r2[12]) );
  DFF_X1 x_r3_reg_12_ ( .D(x_r2[12]), .CK(clk), .Q(x_r3[12]) );
  DFF_X1 x_r1_reg_11_ ( .D(N95), .CK(clk), .Q(x_r1[11]) );
  DFF_X1 x_r2_reg_11_ ( .D(x_r1[11]), .CK(clk), .Q(x_r2[11]) );
  DFF_X1 x_r3_reg_11_ ( .D(x_r2[11]), .CK(clk), .Q(x_r3[11]) );
  DFF_X1 x_r1_reg_10_ ( .D(N96), .CK(clk), .Q(x_r1[10]) );
  DFF_X1 x_r2_reg_10_ ( .D(x_r1[10]), .CK(clk), .Q(x_r2[10]) );
  DFF_X1 x_r3_reg_10_ ( .D(x_r2[10]), .CK(clk), .Q(x_r3[10]) );
  DFF_X1 x_r1_reg_9_ ( .D(N97), .CK(clk), .Q(x_r1[9]) );
  DFF_X1 x_r2_reg_9_ ( .D(x_r1[9]), .CK(clk), .Q(x_r2[9]) );
  DFF_X1 x_r3_reg_9_ ( .D(x_r2[9]), .CK(clk), .Q(x_r3[9]) );
  DFF_X1 x_r1_reg_8_ ( .D(N98), .CK(clk), .Q(x_r1[8]) );
  DFF_X1 x_r2_reg_8_ ( .D(x_r1[8]), .CK(clk), .Q(x_r2[8]) );
  DFF_X1 x_r3_reg_8_ ( .D(x_r2[8]), .CK(clk), .Q(x_r3[8]) );
  DFF_X1 x_r1_reg_7_ ( .D(N99), .CK(clk), .Q(x_r1[7]) );
  DFF_X1 x_r2_reg_7_ ( .D(x_r1[7]), .CK(clk), .Q(x_r2[7]) );
  DFF_X1 x_r3_reg_7_ ( .D(x_r2[7]), .CK(clk), .Q(x_r3[7]) );
  DFF_X1 x_r1_reg_6_ ( .D(N100), .CK(clk), .Q(x_r1[6]) );
  DFF_X1 x_r2_reg_6_ ( .D(x_r1[6]), .CK(clk), .Q(x_r2[6]) );
  DFF_X1 x_r3_reg_6_ ( .D(x_r2[6]), .CK(clk), .Q(x_r3[6]) );
  DFF_X1 x_r1_reg_5_ ( .D(N101), .CK(clk), .Q(x_r1[5]) );
  DFF_X1 x_r2_reg_5_ ( .D(x_r1[5]), .CK(clk), .Q(x_r2[5]) );
  DFF_X1 x_r3_reg_5_ ( .D(x_r2[5]), .CK(clk), .Q(x_r3[5]) );
  DFF_X1 x_r1_reg_4_ ( .D(N102), .CK(clk), .Q(x_r1[4]) );
  DFF_X1 x_r2_reg_4_ ( .D(x_r1[4]), .CK(clk), .Q(x_r2[4]) );
  DFF_X1 x_r3_reg_4_ ( .D(x_r2[4]), .CK(clk), .Q(x_r3[4]) );
  DFF_X1 x_r1_reg_3_ ( .D(N103), .CK(clk), .Q(x_r1[3]) );
  DFF_X1 x_r2_reg_3_ ( .D(x_r1[3]), .CK(clk), .Q(x_r2[3]) );
  DFF_X1 x_r3_reg_3_ ( .D(x_r2[3]), .CK(clk), .Q(x_r3[3]) );
  DFF_X1 x_r1_reg_2_ ( .D(N104), .CK(clk), .Q(x_r1[2]) );
  DFF_X1 x_r2_reg_2_ ( .D(x_r1[2]), .CK(clk), .Q(x_r2[2]) );
  DFF_X1 x_r3_reg_2_ ( .D(x_r2[2]), .CK(clk), .Q(x_r3[2]) );
  DFF_X1 x_r1_reg_1_ ( .D(N105), .CK(clk), .Q(x_r1[1]) );
  DFF_X1 x_r2_reg_1_ ( .D(x_r1[1]), .CK(clk), .Q(x_r2[1]) );
  DFF_X1 x_r3_reg_1_ ( .D(x_r2[1]), .CK(clk), .Q(x_r3[1]) );
  DFF_X1 x_r1_reg_0_ ( .D(N106), .CK(clk), .Q(x_r1[0]) );
  DFF_X1 x_r2_reg_0_ ( .D(x_r1[0]), .CK(clk), .Q(x_r2[0]) );
  DFF_X1 x_r3_reg_0_ ( .D(x_r2[0]), .CK(clk), .Q(x_r3[0]) );
  DFF_X1 x_r4_reg_14_ ( .D(x_r3[14]), .CK(clk), .Q(x_r4[14]) );
  DFF_X1 x_r4_reg_13_ ( .D(x_r3[13]), .CK(clk), .Q(x_r4[13]) );
  DFF_X1 x_r4_reg_12_ ( .D(x_r3[12]), .CK(clk), .Q(x_r4[12]) );
  DFF_X1 x_r4_reg_11_ ( .D(x_r3[11]), .CK(clk), .Q(x_r4[11]) );
  DFF_X1 x_r4_reg_10_ ( .D(x_r3[10]), .CK(clk), .Q(x_r4[10]) );
  DFF_X1 x_r4_reg_9_ ( .D(x_r3[9]), .CK(clk), .Q(x_r4[9]) );
  DFF_X1 x_r4_reg_8_ ( .D(x_r3[8]), .CK(clk), .Q(x_r4[8]) );
  DFF_X1 x_r4_reg_7_ ( .D(x_r3[7]), .CK(clk), .Q(x_r4[7]) );
  DFF_X1 x_r4_reg_6_ ( .D(x_r3[6]), .CK(clk), .Q(x_r4[6]) );
  DFF_X1 x_r4_reg_5_ ( .D(x_r3[5]), .CK(clk), .Q(x_r4[5]) );
  DFF_X1 x_r4_reg_4_ ( .D(x_r3[4]), .CK(clk), .Q(x_r4[4]) );
  DFF_X1 x_r4_reg_3_ ( .D(x_r3[3]), .CK(clk), .Q(x_r4[3]) );
  DFF_X1 x_r4_reg_2_ ( .D(x_r3[2]), .CK(clk), .Q(x_r4[2]) );
  DFF_X1 x_r4_reg_1_ ( .D(x_r3[1]), .CK(clk), .Q(x_r4[1]) );
  DFF_X1 x_r4_reg_0_ ( .D(x_r3[0]), .CK(clk), .Q(x_r4[0]) );
  DFF_X1 c1_r1_reg_17_ ( .D(c1[17]), .CK(clk), .Q(c1_r1[17]) );
  DFF_X1 c1_r1_reg_16_ ( .D(c1[16]), .CK(clk), .Q(c1_r1[16]) );
  DFF_X1 c1_r1_reg_15_ ( .D(c1[15]), .CK(clk), .Q(c1_r1[15]) );
  DFF_X1 c1_r1_reg_14_ ( .D(c1[14]), .CK(clk), .Q(c1_r1[14]) );
  DFF_X1 c1_r1_reg_13_ ( .D(c1[13]), .CK(clk), .Q(c1_r1[13]) );
  DFF_X1 c1_r1_reg_12_ ( .D(c1[12]), .CK(clk), .Q(c1_r1[12]) );
  DFF_X1 c1_r1_reg_11_ ( .D(c1[11]), .CK(clk), .Q(c1_r1[11]) );
  DFF_X1 c1_r1_reg_10_ ( .D(c1[10]), .CK(clk), .Q(c1_r1[10]) );
  DFF_X1 c1_r1_reg_9_ ( .D(c1[9]), .CK(clk), .Q(c1_r1[9]) );
  DFF_X1 c1_r1_reg_8_ ( .D(c1[8]), .CK(clk), .Q(c1_r1[8]) );
  DFF_X1 c1_r1_reg_7_ ( .D(c1[7]), .CK(clk), .Q(c1_r1[7]) );
  DFF_X1 c1_r1_reg_6_ ( .D(c1[6]), .CK(clk), .Q(c1_r1[6]) );
  DFF_X1 c1_r1_reg_5_ ( .D(c1[5]), .CK(clk), .Q(c1_r1[5]) );
  DFF_X1 c1_r1_reg_4_ ( .D(c1[4]), .CK(clk), .Q(c1_r1[4]) );
  DFF_X1 c1_r1_reg_3_ ( .D(c1[3]), .CK(clk), .Q(c1_r1[3]) );
  DFF_X1 c1_r1_reg_2_ ( .D(c1[2]), .CK(clk), .Q(c1_r1[2]) );
  DFF_X1 c1_r1_reg_1_ ( .D(c1[1]), .CK(clk), .Q(c1_r1[1]) );
  DFF_X1 c1_r1_reg_0_ ( .D(c1[0]), .CK(clk), .Q(c1_r1[0]) );
  DFF_X1 c0_r1_reg_17_ ( .D(c0[17]), .CK(clk), .Q(c0_r1[17]) );
  DFF_X1 c0_r2_reg_17_ ( .D(c0_r1[17]), .CK(clk), .Q(c0_r2[17]) );
  DFF_X1 c0_r3_reg_17_ ( .D(c0_r2[17]), .CK(clk), .Q(c0_r3[17]) );
  DFF_X1 c0_r4_reg_17_ ( .D(c0_r3[17]), .CK(clk), .Q(c0_r4[17]) );
  DFF_X1 c0_r1_reg_16_ ( .D(c0[16]), .CK(clk), .Q(c0_r1[16]) );
  DFF_X1 c0_r2_reg_16_ ( .D(c0_r1[16]), .CK(clk), .Q(c0_r2[16]) );
  DFF_X1 c0_r3_reg_16_ ( .D(c0_r2[16]), .CK(clk), .Q(c0_r3[16]) );
  DFF_X1 c0_r4_reg_16_ ( .D(c0_r3[16]), .CK(clk), .Q(c0_r4[16]) );
  DFF_X1 c0_r1_reg_15_ ( .D(c0[15]), .CK(clk), .Q(c0_r1[15]) );
  DFF_X1 c0_r2_reg_15_ ( .D(c0_r1[15]), .CK(clk), .Q(c0_r2[15]) );
  DFF_X1 c0_r3_reg_15_ ( .D(c0_r2[15]), .CK(clk), .Q(c0_r3[15]) );
  DFF_X1 c0_r4_reg_15_ ( .D(c0_r3[15]), .CK(clk), .Q(c0_r4[15]) );
  DFF_X1 c0_r1_reg_14_ ( .D(c0[14]), .CK(clk), .Q(c0_r1[14]) );
  DFF_X1 c0_r2_reg_14_ ( .D(c0_r1[14]), .CK(clk), .Q(c0_r2[14]) );
  DFF_X1 c0_r3_reg_14_ ( .D(c0_r2[14]), .CK(clk), .Q(c0_r3[14]) );
  DFF_X1 c0_r4_reg_14_ ( .D(c0_r3[14]), .CK(clk), .Q(c0_r4[14]) );
  DFF_X1 c0_r1_reg_13_ ( .D(c0[13]), .CK(clk), .Q(c0_r1[13]) );
  DFF_X1 c0_r2_reg_13_ ( .D(c0_r1[13]), .CK(clk), .Q(c0_r2[13]) );
  DFF_X1 c0_r3_reg_13_ ( .D(c0_r2[13]), .CK(clk), .Q(c0_r3[13]) );
  DFF_X1 c0_r4_reg_13_ ( .D(c0_r3[13]), .CK(clk), .Q(c0_r4[13]) );
  DFF_X1 c0_r1_reg_12_ ( .D(c0[12]), .CK(clk), .Q(c0_r1[12]) );
  DFF_X1 c0_r2_reg_12_ ( .D(c0_r1[12]), .CK(clk), .Q(c0_r2[12]) );
  DFF_X1 c0_r3_reg_12_ ( .D(c0_r2[12]), .CK(clk), .Q(c0_r3[12]) );
  DFF_X1 c0_r4_reg_12_ ( .D(c0_r3[12]), .CK(clk), .Q(c0_r4[12]) );
  DFF_X1 c0_r1_reg_11_ ( .D(c0[11]), .CK(clk), .Q(c0_r1[11]) );
  DFF_X1 c0_r2_reg_11_ ( .D(c0_r1[11]), .CK(clk), .Q(c0_r2[11]) );
  DFF_X1 c0_r3_reg_11_ ( .D(c0_r2[11]), .CK(clk), .Q(c0_r3[11]) );
  DFF_X1 c0_r4_reg_11_ ( .D(c0_r3[11]), .CK(clk), .Q(c0_r4[11]) );
  DFF_X1 c0_r1_reg_10_ ( .D(c0[10]), .CK(clk), .Q(c0_r1[10]) );
  DFF_X1 c0_r2_reg_10_ ( .D(c0_r1[10]), .CK(clk), .Q(c0_r2[10]) );
  DFF_X1 c0_r3_reg_10_ ( .D(c0_r2[10]), .CK(clk), .Q(c0_r3[10]) );
  DFF_X1 c0_r4_reg_10_ ( .D(c0_r3[10]), .CK(clk), .Q(c0_r4[10]) );
  DFF_X1 c0_r1_reg_9_ ( .D(c0[9]), .CK(clk), .Q(c0_r1[9]) );
  DFF_X1 c0_r2_reg_9_ ( .D(c0_r1[9]), .CK(clk), .Q(c0_r2[9]) );
  DFF_X1 c0_r3_reg_9_ ( .D(c0_r2[9]), .CK(clk), .Q(c0_r3[9]) );
  DFF_X1 c0_r4_reg_9_ ( .D(c0_r3[9]), .CK(clk), .Q(c0_r4[9]) );
  DFF_X1 c0_r1_reg_8_ ( .D(c0[8]), .CK(clk), .Q(c0_r1[8]) );
  DFF_X1 c0_r2_reg_8_ ( .D(c0_r1[8]), .CK(clk), .Q(c0_r2[8]) );
  DFF_X1 c0_r3_reg_8_ ( .D(c0_r2[8]), .CK(clk), .Q(c0_r3[8]) );
  DFF_X1 c0_r4_reg_8_ ( .D(c0_r3[8]), .CK(clk), .Q(c0_r4[8]) );
  DFF_X1 c0_r1_reg_7_ ( .D(c0[7]), .CK(clk), .Q(c0_r1[7]) );
  DFF_X1 c0_r2_reg_7_ ( .D(c0_r1[7]), .CK(clk), .Q(c0_r2[7]) );
  DFF_X1 c0_r3_reg_7_ ( .D(c0_r2[7]), .CK(clk), .Q(c0_r3[7]) );
  DFF_X1 c0_r4_reg_7_ ( .D(c0_r3[7]), .CK(clk), .Q(c0_r4[7]) );
  DFF_X1 c0_r1_reg_6_ ( .D(c0[6]), .CK(clk), .Q(c0_r1[6]) );
  DFF_X1 c0_r2_reg_6_ ( .D(c0_r1[6]), .CK(clk), .Q(c0_r2[6]) );
  DFF_X1 c0_r3_reg_6_ ( .D(c0_r2[6]), .CK(clk), .Q(c0_r3[6]) );
  DFF_X1 c0_r4_reg_6_ ( .D(c0_r3[6]), .CK(clk), .Q(c0_r4[6]) );
  DFF_X1 c0_r1_reg_5_ ( .D(c0[5]), .CK(clk), .Q(c0_r1[5]) );
  DFF_X1 c0_r2_reg_5_ ( .D(c0_r1[5]), .CK(clk), .Q(c0_r2[5]) );
  DFF_X1 c0_r3_reg_5_ ( .D(c0_r2[5]), .CK(clk), .Q(c0_r3[5]) );
  DFF_X1 c0_r4_reg_5_ ( .D(c0_r3[5]), .CK(clk), .Q(c0_r4[5]) );
  DFF_X1 c0_r1_reg_4_ ( .D(c0[4]), .CK(clk), .Q(c0_r1[4]) );
  DFF_X1 c0_r2_reg_4_ ( .D(c0_r1[4]), .CK(clk), .Q(c0_r2[4]) );
  DFF_X1 c0_r3_reg_4_ ( .D(c0_r2[4]), .CK(clk), .Q(c0_r3[4]) );
  DFF_X1 c0_r4_reg_4_ ( .D(c0_r3[4]), .CK(clk), .Q(c0_r4[4]) );
  DFF_X1 c0_r1_reg_3_ ( .D(c0[3]), .CK(clk), .Q(c0_r1[3]) );
  DFF_X1 c0_r2_reg_3_ ( .D(c0_r1[3]), .CK(clk), .Q(c0_r2[3]) );
  DFF_X1 c0_r3_reg_3_ ( .D(c0_r2[3]), .CK(clk), .Q(c0_r3[3]) );
  DFF_X1 c0_r4_reg_3_ ( .D(c0_r3[3]), .CK(clk), .Q(c0_r4[3]) );
  DFF_X1 c0_r1_reg_2_ ( .D(c0[2]), .CK(clk), .Q(c0_r1[2]) );
  DFF_X1 c0_r2_reg_2_ ( .D(c0_r1[2]), .CK(clk), .Q(c0_r2[2]) );
  DFF_X1 c0_r3_reg_2_ ( .D(c0_r2[2]), .CK(clk), .Q(c0_r3[2]) );
  DFF_X1 c0_r4_reg_2_ ( .D(c0_r3[2]), .CK(clk), .Q(c0_r4[2]) );
  DFF_X1 c0_r1_reg_1_ ( .D(c0[1]), .CK(clk), .Q(c0_r1[1]) );
  DFF_X1 c0_r2_reg_1_ ( .D(c0_r1[1]), .CK(clk), .Q(c0_r2[1]) );
  DFF_X1 c0_r3_reg_1_ ( .D(c0_r2[1]), .CK(clk), .Q(c0_r3[1]) );
  DFF_X1 c0_r4_reg_1_ ( .D(c0_r3[1]), .CK(clk), .Q(c0_r4[1]) );
  DFF_X1 c0_r1_reg_0_ ( .D(c0[0]), .CK(clk), .Q(c0_r1[0]) );
  DFF_X1 c0_r2_reg_0_ ( .D(c0_r1[0]), .CK(clk), .Q(c0_r2[0]) );
  DFF_X1 c0_r3_reg_0_ ( .D(c0_r2[0]), .CK(clk), .Q(c0_r3[0]) );
  DFF_X1 c0_r4_reg_0_ ( .D(c0_r3[0]), .CK(clk), .Q(c0_r4[0]) );
  DFF_X1 c0_r5_reg_17_ ( .D(c0_r4[17]), .CK(clk), .Q(c0_r5[17]) );
  DFF_X1 c0_r5_reg_16_ ( .D(c0_r4[16]), .CK(clk), .Q(c0_r5[16]) );
  DFF_X1 c0_r5_reg_15_ ( .D(c0_r4[15]), .CK(clk), .Q(c0_r5[15]) );
  DFF_X1 c0_r5_reg_14_ ( .D(c0_r4[14]), .CK(clk), .Q(c0_r5[14]) );
  DFF_X1 c0_r5_reg_13_ ( .D(c0_r4[13]), .CK(clk), .Q(c0_r5[13]) );
  DFF_X1 c0_r5_reg_12_ ( .D(c0_r4[12]), .CK(clk), .Q(c0_r5[12]) );
  DFF_X1 c0_r5_reg_11_ ( .D(c0_r4[11]), .CK(clk), .Q(c0_r5[11]) );
  DFF_X1 c0_r5_reg_10_ ( .D(c0_r4[10]), .CK(clk), .Q(c0_r5[10]) );
  DFF_X1 c0_r5_reg_9_ ( .D(c0_r4[9]), .CK(clk), .Q(c0_r5[9]) );
  DFF_X1 c0_r5_reg_8_ ( .D(c0_r4[8]), .CK(clk), .Q(c0_r5[8]) );
  DFF_X1 c0_r5_reg_7_ ( .D(c0_r4[7]), .CK(clk), .Q(c0_r5[7]) );
  DFF_X1 c0_r5_reg_6_ ( .D(c0_r4[6]), .CK(clk), .Q(c0_r5[6]) );
  DFF_X1 c0_r5_reg_5_ ( .D(c0_r4[5]), .CK(clk), .Q(c0_r5[5]) );
  DFF_X1 c0_r5_reg_4_ ( .D(c0_r4[4]), .CK(clk), .Q(c0_r5[4]) );
  DFF_X1 c0_r5_reg_3_ ( .D(c0_r4[3]), .CK(clk), .Q(c0_r5[3]) );
  DFF_X1 c0_r5_reg_2_ ( .D(c0_r4[2]), .CK(clk), .Q(c0_r5[2]) );
  DFF_X1 c0_r5_reg_1_ ( .D(c0_r4[1]), .CK(clk), .Q(c0_r5[1]) );
  DFF_X1 c0_r5_reg_0_ ( .D(c0_r4[0]), .CK(clk), .Q(c0_r5[0]) );
  DFF_X1 sign_r_reg_0_ ( .D(data_in[0]), .CK(clk), .Q(sign_r[0]) );
  DFF_X1 sign_r_reg_1_ ( .D(sign_r[0]), .CK(clk), .Q(sign_r[1]) );
  DFF_X1 sign_r_reg_2_ ( .D(sign_r[1]), .CK(clk), .Q(sign_r[2]) );
  DFF_X1 sign_r_reg_3_ ( .D(sign_r[2]), .CK(clk), .Q(sign_r[3]) );
  DFF_X1 sign_r_reg_4_ ( .D(sign_r[3]), .CK(clk), .Q(sign_r[4]) );
  DFF_X1 sign_r_reg_5_ ( .D(sign_r[4]), .CK(clk), .Q(sign_r[5]) );
  DFF_X1 sign_r_reg_6_ ( .D(sign_r[5]), .CK(clk), .Q(sign_r[6]) );
  DFF_X1 sign_r_reg_7_ ( .D(sign_r[6]), .CK(clk), .Q(sign_r[7]) );
  DFF_X1 sign_r_reg_8_ ( .D(sign_r[7]), .CK(clk), .Q(sign_r[8]), .QN(n12) );
  DFF_X1 valid_in_r_reg_0_ ( .D(N107), .CK(clk), .Q(valid_in_r[0]) );
  DFF_X1 valid_in_r_reg_1_ ( .D(N108), .CK(clk), .Q(valid_in_r[1]) );
  DFF_X1 valid_in_r_reg_2_ ( .D(N109), .CK(clk), .Q(valid_in_r[2]) );
  DFF_X1 valid_in_r_reg_3_ ( .D(N110), .CK(clk), .Q(valid_in_r[3]) );
  DFF_X1 valid_in_r_reg_4_ ( .D(N111), .CK(clk), .Q(valid_in_r[4]) );
  DFF_X1 valid_in_r_reg_5_ ( .D(N112), .CK(clk), .Q(valid_in_r[5]) );
  DFF_X1 valid_in_r_reg_6_ ( .D(N113), .CK(clk), .Q(valid_in_r[6]) );
  DFF_X1 valid_in_r_reg_7_ ( .D(N114), .CK(clk), .Q(valid_in_r[7]) );
  DFF_X1 valid_in_r_reg_8_ ( .D(N115), .CK(clk), .Q(valid_in_r[8]) );
  DFF_X1 sum2_reg_17_ ( .D(N131), .CK(clk), .QN(n58) );
  DFF_X1 sum2_reg_16_ ( .D(N130), .CK(clk), .Q(sum2[16]) );
  DFF_X1 sum2_reg_15_ ( .D(N129), .CK(clk), .Q(sum2[15]) );
  DFF_X1 sum2_reg_14_ ( .D(N128), .CK(clk), .Q(sum2[14]) );
  DFF_X1 sum2_reg_13_ ( .D(N127), .CK(clk), .Q(sum2[13]) );
  DFF_X1 sum2_reg_12_ ( .D(N126), .CK(clk), .Q(sum2[12]) );
  DFF_X1 sum2_reg_11_ ( .D(N125), .CK(clk), .Q(sum2[11]) );
  DFF_X1 sum2_reg_10_ ( .D(N124), .CK(clk), .Q(sum2[10]) );
  DFF_X1 sum2_reg_9_ ( .D(N123), .CK(clk), .Q(sum2[9]) );
  DFF_X1 sum2_reg_8_ ( .D(N122), .CK(clk), .Q(sum2[8]) );
  DFF_X1 sum2_reg_7_ ( .D(N121), .CK(clk), .Q(sum2[7]) );
  DFF_X1 sum2_reg_6_ ( .D(N120), .CK(clk), .Q(sum2[6]) );
  DFF_X1 sum2_reg_5_ ( .D(N119), .CK(clk), .Q(sum2[5]) );
  DFF_X1 sum2_reg_4_ ( .D(N118), .CK(clk), .Q(sum2[4]) );
  DFF_X1 sum2_reg_3_ ( .D(N117), .CK(clk), .Q(sum2[3]) );
  DFF_X1 sum2_reg_2_ ( .D(N116), .CK(clk), .Q(sum2[2]) );
  DFF_X1 sum2_rnd_reg_14_ ( .D(n57), .CK(clk), .QN(n29) );
  DFF_X1 sum2_rnd_reg_13_ ( .D(n28), .CK(clk), .QN(n30) );
  DFF_X1 sum2_rnd_reg_12_ ( .D(n27), .CK(clk), .QN(n31) );
  DFF_X1 sum2_rnd_reg_11_ ( .D(n26), .CK(clk), .QN(n32) );
  DFF_X1 sum2_rnd_reg_10_ ( .D(n25), .CK(clk), .QN(n33) );
  DFF_X1 sum2_rnd_reg_9_ ( .D(n24), .CK(clk), .QN(n34) );
  DFF_X1 sum2_rnd_reg_8_ ( .D(n23), .CK(clk), .QN(n35) );
  DFF_X1 sum2_rnd_reg_7_ ( .D(n22), .CK(clk), .QN(n36) );
  DFF_X1 sum2_rnd_reg_6_ ( .D(n1), .CK(clk), .QN(n37) );
  DFF_X1 sum2_rnd_reg_5_ ( .D(n940), .CK(clk), .QN(n38) );
  DFF_X1 sum2_rnd_reg_4_ ( .D(n930), .CK(clk), .QN(n39) );
  DFF_X1 sum2_rnd_reg_3_ ( .D(n920), .CK(clk), .QN(n40) );
  DFF_X1 sum2_rnd_reg_2_ ( .D(n911), .CK(clk), .QN(n41) );
  DFF_X1 sum2_rnd_reg_1_ ( .D(n900), .CK(clk), .QN(n42) );
  DFF_X1 sum2_rnd_reg_0_ ( .D(n890), .CK(clk), .QN(n43) );
  DFF_X1 valid_out_reg ( .D(N147), .CK(clk), .Q(valid_out) );
  DFF_X1 data_out_reg_15_ ( .D(N197), .CK(clk), .Q(data_out[15]) );
  DFF_X1 data_out_reg_14_ ( .D(N196), .CK(clk), .Q(data_out[14]) );
  DFF_X1 data_out_reg_13_ ( .D(N195), .CK(clk), .Q(data_out[13]) );
  DFF_X1 data_out_reg_12_ ( .D(N194), .CK(clk), .Q(data_out[12]) );
  DFF_X1 data_out_reg_11_ ( .D(N193), .CK(clk), .Q(data_out[11]) );
  DFF_X1 data_out_reg_10_ ( .D(N192), .CK(clk), .Q(data_out[10]) );
  DFF_X1 data_out_reg_9_ ( .D(N191), .CK(clk), .Q(data_out[9]) );
  DFF_X1 data_out_reg_8_ ( .D(N190), .CK(clk), .Q(data_out[8]) );
  DFF_X1 data_out_reg_7_ ( .D(N189), .CK(clk), .Q(data_out[7]) );
  DFF_X1 data_out_reg_6_ ( .D(N188), .CK(clk), .Q(data_out[6]) );
  DFF_X1 data_out_reg_5_ ( .D(N187), .CK(clk), .Q(data_out[5]) );
  DFF_X1 data_out_reg_4_ ( .D(N186), .CK(clk), .Q(data_out[4]) );
  DFF_X1 data_out_reg_3_ ( .D(N185), .CK(clk), .Q(data_out[3]) );
  DFF_X1 data_out_reg_2_ ( .D(N184), .CK(clk), .Q(data_out[2]) );
  DFF_X1 data_out_reg_1_ ( .D(N183), .CK(clk), .Q(data_out[1]) );
  DFF_X1 data_out_reg_0_ ( .D(N182), .CK(clk), .Q(data_out[0]) );
  gng_lzd u_gng_lzd ( .data_in(data_in[63:3]), .data_out(num_lzd) );
  gng_coef u_gng_coef ( .clk(clk), .addr({num_lzd_r, offset}), .c0(c0), .c1(c1), .c2(c2) );
  gng_smul_16_18_sadd_37 u_gng_smul_16_18_sadd_37 ( .clk(clk), .a({1'b0, x_r1}), .b({1'b0, c2}), .c({c1_r1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .p({sum1, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20}) );
  gng_smul_16_18 u_gng_smul_16_18 ( .clk(clk), .a({1'b0, x_r4}), .b(sum1), .p(
        {SYNOPSYS_UNCONNECTED_21, mul1, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40}) );
  gng_interp_DW01_inc_0 add_219 ( .A({1'b1, n29, n30, n31, n32, n33, n34, n35, 
        n36, n37, n38, n39, n40, n41, n42, n43}), .SUM({N181, N180, N179, N178, 
        N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, 
        SYNOPSYS_UNCONNECTED_41}) );
  gng_interp_DW01_add_1 add_199 ( .A(c0_r5), .B({mul1[32], mul1[32], mul1[32], 
        mul1[32], mul1}), .CI(1'b0), .SUM({N131, N130, N129, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43}) );
  NOR2_X1 U3 ( .A1(n980), .A2(n55), .ZN(N197) );
  INV_X1 U4 ( .A(N181), .ZN(n980) );
  NAND2_X1 U5 ( .A1(n49), .A2(n47), .ZN(N71) );
  NAND2_X1 U6 ( .A1(n48), .A2(n47), .ZN(N72) );
  NAND2_X1 U8 ( .A1(n46), .A2(n47), .ZN(N73) );
  NAND2_X1 U9 ( .A1(n52), .A2(n45), .ZN(N62) );
  NAND2_X1 U10 ( .A1(n51), .A2(n45), .ZN(N66) );
  NAND2_X1 U11 ( .A1(n47), .A2(n45), .ZN(N70) );
  NAND2_X1 U12 ( .A1(n51), .A2(n49), .ZN(N67) );
  NAND2_X1 U13 ( .A1(n51), .A2(n48), .ZN(N68) );
  NAND2_X1 U14 ( .A1(n51), .A2(n46), .ZN(N69) );
  NAND2_X1 U15 ( .A1(n52), .A2(n49), .ZN(N63) );
  NAND2_X1 U16 ( .A1(n52), .A2(n48), .ZN(N64) );
  NAND2_X1 U17 ( .A1(n52), .A2(n46), .ZN(N65) );
  AND2_X1 U18 ( .A1(num_lzd[0]), .A2(n970), .ZN(N6) );
  AND2_X1 U19 ( .A1(num_lzd[1]), .A2(n970), .ZN(N7) );
  AND2_X1 U20 ( .A1(num_lzd[3]), .A2(n960), .ZN(N9) );
  AND2_X1 U21 ( .A1(num_lzd[2]), .A2(n960), .ZN(N8) );
  AND2_X1 U22 ( .A1(num_lzd[4]), .A2(n960), .ZN(N10) );
  AND2_X1 U23 ( .A1(num_lzd[5]), .A2(n970), .ZN(N11) );
  NAND2_X1 U24 ( .A1(sign_r[8]), .A2(n960), .ZN(n55) );
  NAND2_X1 U25 ( .A1(n960), .A2(n12), .ZN(n56) );
  BUF_X1 U26 ( .A(rstn), .Z(n960) );
  BUF_X1 U27 ( .A(rstn), .Z(n970) );
  OAI22_X1 U28 ( .A1(n55), .A2(n43), .B1(n43), .B2(n56), .ZN(N182) );
  OAI22_X1 U29 ( .A1(n55), .A2(n1120), .B1(n42), .B2(n56), .ZN(N183) );
  INV_X1 U30 ( .A(N167), .ZN(n1120) );
  OAI22_X1 U31 ( .A1(n55), .A2(n1111), .B1(n41), .B2(n56), .ZN(N184) );
  INV_X1 U32 ( .A(N168), .ZN(n1111) );
  OAI22_X1 U33 ( .A1(n55), .A2(n1100), .B1(n40), .B2(n56), .ZN(N185) );
  INV_X1 U34 ( .A(N169), .ZN(n1100) );
  OAI22_X1 U35 ( .A1(n55), .A2(n1090), .B1(n39), .B2(n56), .ZN(N186) );
  INV_X1 U36 ( .A(N170), .ZN(n1090) );
  OAI22_X1 U37 ( .A1(n55), .A2(n1080), .B1(n38), .B2(n56), .ZN(N187) );
  INV_X1 U38 ( .A(N171), .ZN(n1080) );
  OAI22_X1 U39 ( .A1(n55), .A2(n1070), .B1(n37), .B2(n56), .ZN(N188) );
  INV_X1 U40 ( .A(N172), .ZN(n1070) );
  OAI22_X1 U41 ( .A1(n55), .A2(n1060), .B1(n36), .B2(n56), .ZN(N189) );
  INV_X1 U42 ( .A(N173), .ZN(n1060) );
  OAI22_X1 U43 ( .A1(n55), .A2(n1050), .B1(n35), .B2(n56), .ZN(N190) );
  INV_X1 U44 ( .A(N174), .ZN(n1050) );
  OAI22_X1 U45 ( .A1(n55), .A2(n1040), .B1(n34), .B2(n56), .ZN(N191) );
  INV_X1 U46 ( .A(N175), .ZN(n1040) );
  OAI22_X1 U47 ( .A1(n55), .A2(n1030), .B1(n33), .B2(n56), .ZN(N192) );
  INV_X1 U48 ( .A(N176), .ZN(n1030) );
  OAI22_X1 U49 ( .A1(n55), .A2(n1020), .B1(n32), .B2(n56), .ZN(N193) );
  INV_X1 U50 ( .A(N177), .ZN(n1020) );
  OAI22_X1 U51 ( .A1(n55), .A2(n1011), .B1(n31), .B2(n56), .ZN(N194) );
  INV_X1 U52 ( .A(N178), .ZN(n1011) );
  OAI22_X1 U53 ( .A1(n55), .A2(n1000), .B1(n30), .B2(n56), .ZN(N195) );
  INV_X1 U54 ( .A(N179), .ZN(n1000) );
  OAI22_X1 U55 ( .A1(n55), .A2(n990), .B1(n29), .B2(n56), .ZN(N196) );
  INV_X1 U56 ( .A(N180), .ZN(n990) );
  AND3_X1 U57 ( .A1(n44), .A2(n810), .A3(num_lzd_r[2]), .ZN(n51) );
  AND2_X1 U58 ( .A1(n50), .A2(num_lzd_r[3]), .ZN(n47) );
  AND2_X1 U59 ( .A1(n50), .A2(n810), .ZN(n52) );
  NAND4_X1 U60 ( .A1(num_lzd_r[3]), .A2(num_lzd_r[2]), .A3(n44), .A4(n45), 
        .ZN(N74) );
  AND3_X1 U61 ( .A1(num_lzd_r[4]), .A2(n970), .A3(num_lzd_r[5]), .ZN(n44) );
  AND4_X1 U62 ( .A1(n960), .A2(n710), .A3(num_lzd_r[5]), .A4(n54), .ZN(n53) );
  NOR3_X1 U63 ( .A1(n1010), .A2(n910), .A3(n810), .ZN(n54) );
  NAND2_X1 U64 ( .A1(n53), .A2(num_lzd_r[0]), .ZN(N61) );
  AND2_X1 U65 ( .A1(n44), .A2(n910), .ZN(n50) );
  NAND2_X1 U66 ( .A1(n53), .A2(n1110), .ZN(N60) );
  AND2_X1 U67 ( .A1(data_in[6]), .A2(n960), .ZN(N88) );
  AND2_X1 U68 ( .A1(data_in[14]), .A2(n960), .ZN(N80) );
  AND2_X1 U69 ( .A1(data_in[10]), .A2(n970), .ZN(N84) );
  AND2_X1 U70 ( .A1(n970), .A2(data_in[3]), .ZN(N91) );
  AND2_X1 U71 ( .A1(data_in[16]), .A2(n960), .ZN(N78) );
  AND2_X1 U72 ( .A1(data_in[15]), .A2(n960), .ZN(N79) );
  AND2_X1 U73 ( .A1(data_in[13]), .A2(n960), .ZN(N81) );
  AND2_X1 U74 ( .A1(data_in[12]), .A2(n960), .ZN(N82) );
  AND2_X1 U75 ( .A1(data_in[11]), .A2(n960), .ZN(N83) );
  AND2_X1 U76 ( .A1(data_in[9]), .A2(n960), .ZN(N85) );
  AND2_X1 U77 ( .A1(data_in[8]), .A2(n960), .ZN(N86) );
  AND2_X1 U78 ( .A1(data_in[7]), .A2(n960), .ZN(N87) );
  AND2_X1 U79 ( .A1(data_in[5]), .A2(n960), .ZN(N89) );
  AND2_X1 U80 ( .A1(data_in[4]), .A2(n960), .ZN(N90) );
  AND2_X1 U81 ( .A1(valid_in_r[8]), .A2(n970), .ZN(N147) );
  AND2_X1 U82 ( .A1(valid_in_r[7]), .A2(n970), .ZN(N115) );
  AND2_X1 U83 ( .A1(valid_in_r[6]), .A2(n970), .ZN(N114) );
  AND2_X1 U84 ( .A1(valid_in_r[5]), .A2(n970), .ZN(N113) );
  AND2_X1 U85 ( .A1(valid_in_r[4]), .A2(n970), .ZN(N112) );
  AND2_X1 U86 ( .A1(valid_in_r[3]), .A2(n970), .ZN(N111) );
  AND2_X1 U87 ( .A1(valid_in_r[2]), .A2(n970), .ZN(N110) );
  AND2_X1 U88 ( .A1(valid_in_r[1]), .A2(n970), .ZN(N109) );
  AND2_X1 U89 ( .A1(valid_in_r[0]), .A2(n970), .ZN(N108) );
  AND2_X1 U90 ( .A1(valid_in), .A2(n970), .ZN(N107) );
  AND2_X1 U91 ( .A1(data_in[17]), .A2(n970), .ZN(N77) );
  AND2_X1 U92 ( .A1(data_in[2]), .A2(n970), .ZN(N75) );
  AND2_X1 U93 ( .A1(data_in[1]), .A2(n970), .ZN(N76) );
  XOR2_X1 U94 ( .A(sum2[9]), .B(n610), .Z(n1) );
  AND2_X1 U95 ( .A1(sum2[2]), .A2(sum2[3]), .ZN(n3) );
  AND2_X1 U96 ( .A1(sum2[4]), .A2(n3), .ZN(n4) );
  AND2_X1 U97 ( .A1(sum2[7]), .A2(n17), .ZN(n5) );
  AND2_X1 U98 ( .A1(sum2[8]), .A2(n5), .ZN(n610) );
  AND2_X1 U99 ( .A1(sum2[9]), .A2(n610), .ZN(n13) );
  AND2_X1 U100 ( .A1(sum2[12]), .A2(n19), .ZN(n14) );
  AND2_X1 U101 ( .A1(sum2[15]), .A2(n21), .ZN(n15) );
  AND2_X1 U102 ( .A1(sum2[5]), .A2(n4), .ZN(n16) );
  AND2_X1 U103 ( .A1(sum2[6]), .A2(n16), .ZN(n17) );
  AND2_X1 U104 ( .A1(sum2[10]), .A2(n13), .ZN(n18) );
  AND2_X1 U105 ( .A1(sum2[11]), .A2(n18), .ZN(n19) );
  AND2_X1 U106 ( .A1(sum2[13]), .A2(n14), .ZN(n20) );
  AND2_X1 U107 ( .A1(sum2[14]), .A2(n20), .ZN(n21) );
  XOR2_X1 U108 ( .A(sum2[10]), .B(n13), .Z(n22) );
  XOR2_X1 U109 ( .A(sum2[11]), .B(n18), .Z(n23) );
  XOR2_X1 U110 ( .A(sum2[12]), .B(n19), .Z(n24) );
  XOR2_X1 U111 ( .A(sum2[13]), .B(n14), .Z(n25) );
  XOR2_X1 U112 ( .A(sum2[14]), .B(n20), .Z(n26) );
  XOR2_X1 U113 ( .A(sum2[15]), .B(n21), .Z(n27) );
  XOR2_X1 U114 ( .A(sum2[16]), .B(n15), .Z(n28) );
  XOR2_X1 U115 ( .A(n58), .B(n950), .Z(n57) );
  NAND2_X1 U116 ( .A1(sum2[16]), .A2(n15), .ZN(n950) );
  NOR2_X1 U117 ( .A1(num_lzd_r[1]), .A2(num_lzd_r[0]), .ZN(n45) );
  NOR2_X1 U118 ( .A1(n1110), .A2(num_lzd_r[1]), .ZN(n49) );
  NOR2_X1 U119 ( .A1(n1010), .A2(num_lzd_r[0]), .ZN(n48) );
  NOR2_X1 U120 ( .A1(n1010), .A2(n1110), .ZN(n46) );
  NOR2_X1 U121 ( .A1(n59), .A2(n600), .ZN(N106) );
  NOR2_X1 U122 ( .A1(n611), .A2(n620), .ZN(N105) );
  NOR2_X1 U123 ( .A1(n630), .A2(n640), .ZN(N104) );
  NOR2_X1 U124 ( .A1(n650), .A2(n660), .ZN(N103) );
  NOR2_X1 U125 ( .A1(n670), .A2(n680), .ZN(N102) );
  NOR2_X1 U126 ( .A1(n690), .A2(n700), .ZN(N101) );
  NOR2_X1 U127 ( .A1(n711), .A2(n720), .ZN(N100) );
  NOR2_X1 U128 ( .A1(n730), .A2(n740), .ZN(N99) );
  NOR2_X1 U129 ( .A1(n750), .A2(n760), .ZN(N98) );
  NOR2_X1 U130 ( .A1(n770), .A2(n780), .ZN(N97) );
  NOR2_X1 U131 ( .A1(n790), .A2(n800), .ZN(N96) );
  NOR2_X1 U132 ( .A1(n811), .A2(n820), .ZN(N95) );
  NOR2_X1 U133 ( .A1(n830), .A2(n840), .ZN(N94) );
  NOR2_X1 U134 ( .A1(n850), .A2(n860), .ZN(N93) );
  NOR2_X1 U135 ( .A1(n870), .A2(n880), .ZN(N92) );
  XOR2_X1 U136 ( .A(sum2[2]), .B(sum2[3]), .Z(n890) );
  XOR2_X1 U137 ( .A(sum2[4]), .B(n3), .Z(n900) );
  XOR2_X1 U138 ( .A(sum2[5]), .B(n4), .Z(n911) );
  XOR2_X1 U139 ( .A(sum2[6]), .B(n16), .Z(n920) );
  XOR2_X1 U140 ( .A(sum2[7]), .B(n17), .Z(n930) );
  XOR2_X1 U141 ( .A(sum2[8]), .B(n5), .Z(n940) );
endmodule


module gng ( clk, rstn, ce, valid_out, data_out );
  output [15:0] data_out;
  input clk, rstn, ce;
  output valid_out;
  wire   valid_out_ctg;
  wire   [63:0] data_out_ctg;

  gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff u_gng_ctg ( .clk(
        clk), .rstn(rstn), .ce(ce), .valid_out(valid_out_ctg), .data_out(
        data_out_ctg) );
  gng_interp u_gng_interp ( .clk(clk), .rstn(rstn), .valid_in(valid_out_ctg), 
        .data_in(data_out_ctg), .valid_out(valid_out), .data_out(data_out) );
endmodule

