* Nettran: AMD.64 Release B-2008.09.SP5.26004 2012/07/19
* Created:  4/21/2018  16:00
* Options: -rootCell gng -verilog-b0 VSS -verilog-b1 VDD -sp /home/standard_cell_libraries/NangateOpenCellLibrary_PDKv1_3_v2010_12/lib/Back_End/spice/NangateOpenCellLibrary.spi -verilog /home/mohamed/Desktop/ref_flow/pnr/output_verilog_withphysical -outType spice -outName gng.sp 

.GLOBAL VDD VSS 

.SUBCKT XOR2_X2 A B Z VDD VSS 
M_i_41_29 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47_27 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_18 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_35 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19_23 net_001b A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24_4 VSS B net_001b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XNOR2_X2 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_25 VDD B net_003b VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48_8 net_003b A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42_14 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_23_12 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17_20 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11_23 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT TLAT_X1 D G OE Q VDD VSS 
M_i_111 Q net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_106 net_010 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_91 net_005 OE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_99 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 VDD net_006 net_009 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_81 net_009 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_003 net_000 net_008 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_70 net_008 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_64 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 Q OE net_007 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_47 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_34 net_005 OE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TINV_X1 EN I ZN VDD VSS 
M_i_29 ZN EN net_002 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24 net_002 I VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VDD EN net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 ZN net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_7 net_001 I VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0 VSS EN net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TBUF_X8 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X4 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X2 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X16 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_10 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_83 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_42 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_51 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9_17 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18_103 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39_66 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50_12 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_116 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_106 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_120 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_43 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42_108 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37_112 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45_122 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40_125 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X1 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT SDFF_X2 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_115_2 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108_51 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7_4 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_50 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFF_X1 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFS_X2 D SE SI SN CK Q QN VDD VSS 
M_i_230_17 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237_1 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103_26 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110_2 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 VSS net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_93 net_014 SN net_015 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFS_X1 D SE SI SN CK Q QN VDD VSS 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 net_015 net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_93 net_014 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFR_X2 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_116_1 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123_146 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_10 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7_145 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFR_X1 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X2 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_277_67 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290_11 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 net_013 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_106 net_017 SN net_016 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_119 net_019 RN net_018 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_114 net_018 net_017 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_125_68 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132_2 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X1 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_106 net_017 net_013 net_016 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_114 net_018 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_119 net_019 net_017 net_018 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 ZN_neg A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT OR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_1__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m0 VDD A2 net_0__m0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m0 net_0__m0_0__m0_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m1 ZN_neg A1 net_0__m0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m1 net_0__m0_0__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 ZN VDD VSS 
M_i_8 VDD A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 B3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 ZN A3 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_0 B3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 VDD A2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_1__m3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN A1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_1__m2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 VDD B2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 net_2__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN B1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 net_2__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_1 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_0 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_5 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 A1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_0 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_1 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_5 A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 ZN A1 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A2 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 ZN C1 net_4__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 net_4__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 VDD C2 net_4__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 net_4__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0__m1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_3_x4_0 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_1 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_2 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_3 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN_4 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_4 C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_7_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 VDD B2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 net_1__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN B1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_1__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X4 A B C1 C2 ZN VDD VSS 
M_i_5__m3 VDD C2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_2__m3 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN C1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_2__m2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_0 A net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_1__m3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7_1_96 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_102 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34_44 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_56 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_88 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24_95 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_68 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6_75 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8_108 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_109 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_8 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29_45 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_52 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_79 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13_89 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_77 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22_71 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5_83 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_65 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_56 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_52 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_43 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_34 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_24 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_85 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_67 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_58 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_49 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_40 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_31 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5_1_m2__m1 VDD A3 net_1_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m1 net_1_0__m1 A2 net_0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m1 net_0_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m0 ZN A1 net_0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m0 net_0_0__m0_0 A2 net_1_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1_m2__m0 net_1_0__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0_x2__m1 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m1 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m0 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2__m0 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_52 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_154 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_49 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_100 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_202 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_87 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_36 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_189 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_15 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_66 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_168 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_17 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_68 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_170 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_43 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_94 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_196 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_75 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_24 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_177 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_34 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_85 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_187 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5__m3 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m3 VSS A3 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m3 net_1__m3 A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5__m0_x2__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_2__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_x2__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m1 VSS A2 net_0__m0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X2 A B S Z VDD VSS 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_1_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 Z_neg B net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_2 x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS x1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT LOGIC1_X1 Z VDD VSS 
M_p_tran_2 VDD A Z VDD PMOS_VTL L=0.050000U W=0.135000U 
M_n_tran_1 VSS A A VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT FILLCELL_X1 VDD VSS 
.ENDS

.SUBCKT DLL_X2 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_92_11 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_42_3 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLL_X1 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X2 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_89 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_41 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X1 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X2 D SN CK Q QN VDD VSS 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189_10 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182_20 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86_15 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79_29 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X1 D SN CK Q QN VDD VSS 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X2 D RN CK Q QN VDD VSS 
M_i_187_39 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180_3 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83_49 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76_4 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X1 D RN CK Q QN VDD VSS 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFRS_X2 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP81_1_55 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0_51 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 z41 z56 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN51 VSS RN nn5 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN91_0_0_58 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81_53 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFFRS_X1 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 RN z56 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN51 VSS z41 nn5 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X8 CK E GCK VDD VSS 
M_i_109_4_19_36 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24_52 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_22 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_53 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74_97 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71_87 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_99 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_72 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57_165 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7_25_30 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10_28 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_58 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_40 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66_78 VSS net_000 net_007d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75_82 net_007d CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_71 net_007c CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_63 VSS net_000 net_007c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_174 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X4 CK E GCK VDD VSS 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X2 CK E GCK VDD VSS 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X1 CK E GCK VDD VSS 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X8 CK E SE GCK VDD VSS 
M_i_133_10_28_7 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11_14 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_20 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_38 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72_145 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69_164 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_158 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_163 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101_94 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29_4 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15_27 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_55 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_12 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76_137 net_008d CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77_169 net_007 net_002 net_008d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_123 net_007 net_002 net_008c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_150 net_008c CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33_93 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X4 CK E SE GCK VDD VSS 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X2 CK E SE GCK VDD VSS 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X1 CK E SE GCK VDD VSS 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT BUF_X8 A Z VDD VSS 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X4 A Z VDD VSS 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 VSS B2 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_1__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 ZN B1 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 net_1__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_0 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_1 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A2 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_5 A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_1 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_0 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 C1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_5 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_7__m0 net_3 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0 net_0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_2__m0_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN C1 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_2__m1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_0_x4_3 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_2 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_1 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_0 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN_4 C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_4 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 net_2 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS B2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN B1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS B2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN B1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m0_x2__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m0 VSS B2 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 net_0__m0_0__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 ZN B1 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_0__m0_0__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X4 A B C1 C2 ZN VDD VSS 
M_i_11_3 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_2 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_0 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_1 VDD ZN_3 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_0 ZN_4 ZN_3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 C2 ZN_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_3 C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10_3 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_2 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_1 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_1 VSS ZN_3 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_0 ZN_4 ZN_3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 net_1 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1 B net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT ANTENNA_X1 A VDD VSS 
.ENDS

.SUBCKT AND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 x1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A2 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 x1 A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A1 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 x1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 VDD A3 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 x1 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0__m1 A1 x1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 x1 A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_0_x4_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m1 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m0 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_4__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 VSS A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT FILLCELL_X2 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X4 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X8 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X16 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X32 VDD VSS 
.ENDS

.SUBCKT NAND2_X4 A1 A2 ZN VDD VSS 
M_i_2_3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_3 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_2 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_0 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X4 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m1_58 VDD A2 net_0__m0__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1_45 net_0__m0__m2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0_52 ZN A1 net_0__m0__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0_38 net_0__m0__m3 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m1_23 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1_57 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0_35 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0_16 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFF_X2 D CK Q QN VDD VSS 
M_MP13_26 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14_5 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13_38 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14_8 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKBUF_X3 A Z VDD VSS 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN C1 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_2 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 ZN C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NOR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X2 A Z VDD VSS 
M_i_1_0_x2_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X1 A B S Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B net_3 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_3 x1 Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_5 Z_neg x1 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_1 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 VDD A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X16 A Z VDD VSS 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X2 A ZN VDD VSS 
M_i_1_0_x2_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT LOGIC0_X1 Z VDD VSS 
M_transistor_0 VDD A A VDD PMOS_VTL L=0.050000U W=0.090000U 
M_n_tran_1 VSS A Z VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT DFF_X1 D CK Q QN VDD VSS 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKBUF_X2 A Z VDD VSS 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT XNOR2_X1 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NOR2_X1 A1 A2 ZN VDD VSS 
M_i_2 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X1 A1 A2 ZN VDD VSS 
M_i_2 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XOR2_X1 A B Z VDD VSS 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AND2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT INV_X4 A ZN VDD VSS 
M_i_1_0_x4_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X8 A ZN VDD VSS 
M_i_1_0_x8_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x8_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X32 A Z VDD VSS 
M_i_1_31 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_14 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_13 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_12 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_11 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_10 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_9 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_15 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_14 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_13 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_12 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_11 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_10 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_9 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_8 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT HA_X1 A B CO S VDD VSS 
M_i_11 CO CO_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15 VDD B CO_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_14 CO_neg A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 x1 A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_2 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD x1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 A S VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 S B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 CO CO_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS B net_3 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_12 net_3 A CO_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_6 VSS A x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 x1 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS x1 S VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 S A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VSS B net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X1 A ZN VDD VSS 
M_i_1 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT FA_X1 A B CI CO S VDD VSS 
M_instance_315 S net_005 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_275 VDD A net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_280 net_009 B net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_284 net_010 CI net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_290 net_005 net_001 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_303 net_011 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_297 VDD CI net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_309 net_011 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_263 VDD B net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_269 net_008 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_257 net_001 CI net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_251 net_007 A net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_246 VDD B net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_239 CO net_001 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_233 S net_005 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_instance_194 VSS A net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_199 net_003 B net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_203 net_004 CI net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_209 net_005 net_001 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_221 net_006 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_215 VSS CI net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_227 net_006 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_182 VSS B net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_188 net_002 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_176 net_001 CI net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_170 net_000 A net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_166 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_159 CO net_001 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X16 A ZN VDD VSS 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKBUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.095000U 
.ENDS

.SUBCKT BUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT INV_X32 A ZN VDD VSS 
M_i_1_31 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT gng_lzd data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] 
+ VDD VSS data_in[60] data_in[59] data_in[58] data_in[57] data_in[56] data_in[55] 
+ data_in[54] data_in[53] data_in[52] data_in[51] data_in[50] data_in[49] data_in[48] 
+ data_in[47] data_in[46] data_in[45] data_in[44] data_in[43] data_in[42] data_in[41] 
+ data_in[40] data_in[39] data_in[38] data_in[37] data_in[36] data_in[35] data_in[34] 
+ data_in[33] data_in[32] data_in[31] data_in[30] data_in[29] data_in[28] data_in[27] 
+ data_in[26] data_in[25] data_in[24] data_in[23] data_in[22] data_in[21] data_in[20] 
+ data_in[19] data_in[18] data_in[17] data_in[16] data_in[15] data_in[14] data_in[13] 
+ data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] data_in[7] data_in[6] 
+ data_in[5] data_in[4] data_in[3] data_in[2] data_in[1] data_in[0] 
XU22 n58 n15 n18 n14 n56 VDD VSS OAI22_X1 
XU21 n54 n34 n33 n39 n51 VDD VSS OAI22_X1 
XU20 n45 n5 VDD VSS INV_X1 
XU19 n48 n22 VDD VSS INV_X1 
XU18 data_out[5] n48 n43 VDD VSS NAND2_X1 
XU17 n55 n2 VDD VSS INV_X1 
XU16 n55 n130 n42 VDD VSS NAND2_X1 
XU15 n42 n43 data_out[4] VDD VSS NAND2_X1 
XU14 n55 n56 n57 n2 n49 VDD VSS AOI22_X1 
XU13 n48 n51 n52 n22 n50 VDD VSS AOI22_X1 
XU12 data_out[5] n49 n50 n130 n134 VDD VSS OAI22_X1 
XU11 n130 n48 n24 n46 VDD VSS NOR3_X1 
XU10 n46 n45 n2 n44 VDD VSS AOI21_X1 
XU9 n44 n33 n43 n14 n42 n131 VDD VSS OAI221_X1 
XU8 n55 n70 n71 n2 n59 VDD VSS AOI22_X1 
XU7 n67 n37 n68 n35 n69 n40 n60 VDD VSS AOI222_X1 
XU6 n61 data_out[5] n59 n60 n43 n133 VDD VSS OAI221_X1 
XU5 n91 n92 n93 n94 n83 VDD VSS NOR4_X1 
XU4 n85 n86 n87 n88 n84 VDD VSS NOR4_X1 
XU3 n82 n130 n55 n83 n84 n42 n132 VDD VSS OAI222_X1 
XU2 data_in[55] data_in[56] data_in[54] n98 n45 VDD VSS NOR4_X1 
XU76 data_in[13] n23 data_in[15] data_in[14] n48 VDD VSS NOR4_X1 
XU44 data_in[45] n4 data_in[47] data_in[46] n55 VDD VSS NOR4_X2 
XU117 data_in[47] n11 VDD VSS INV_X1 
XU116 data_in[35] n19 VDD VSS INV_X1 
XU115 data_in[51] n10 VDD VSS INV_X1 
XU114 n89 data_in[44] n78 VDD VSS OR2_X1 
XU113 n95 data_in[60] n73 VDD VSS OR2_X1 
XU112 data_in[26] n27 VDD VSS INV_X1 
XU111 n64 data_in[27] n27 n102 VDD VSS OAI21_X1 
XU110 data_in[43] n16 VDD VSS INV_X1 
XU109 n78 data_in[42] n16 n88 VDD VSS AOI21_X1 
XU108 data_in[59] n7 VDD VSS INV_X1 
XU107 n73 data_in[58] n7 n94 VDD VSS AOI21_X1 
XU106 n114 data_in[12] n68 VDD VSS NOR2_X1 
XU105 n108 data_in[28] n64 VDD VSS NOR2_X1 
XU104 data_in[2] data_in[1] data_in[4] data_in[3] n113 VDD VSS NOR4_X1 
XU103 data_in[37] n15 n99 VDD VSS OR2_X1 
XU102 data_in[39] data_in[40] data_in[38] n99 n58 VDD VSS NOR4_X1 
XU101 data_in[23] n28 VDD VSS INV_X1 
XU100 data_in[27] n26 VDD VSS INV_X1 
XU99 n65 n28 n63 n26 n64 n62 VDD VSS AOI221_X1 
XU98 n62 n48 n130 n61 VDD VSS OR3_X1 
XU97 data_in[0] n33 n39 n112 VDD VSS OR3_X1 
XU96 n58 data_in[40] n15 n77 VDD VSS OR3_X1 
XU95 n45 data_in[56] n6 n72 VDD VSS OR3_X1 
XU94 data_in[6] n38 VDD VSS INV_X1 
XU93 n67 data_in[7] n38 n109 VDD VSS OAI21_X1 
XU92 data_in[22] n29 VDD VSS INV_X1 
XU91 n63 data_in[23] n29 n103 VDD VSS OAI21_X1 
XU90 data_in[2] n41 VDD VSS INV_X1 
XU89 n69 data_in[3] n41 n110 VDD VSS OAI21_X1 
XU88 data_in[18] n31 VDD VSS INV_X1 
XU87 n66 data_in[19] n31 n104 VDD VSS OAI21_X1 
XU86 data_in[14] n32 VDD VSS INV_X1 
XU85 n106 data_in[15] n32 n105 VDD VSS OAI21_X1 
XU84 n80 n13 VDD VSS INV_X1 
XU83 n13 data_in[30] n20 n85 VDD VSS AOI21_X1 
XU82 n4 data_in[46] n11 n91 VDD VSS AOI21_X1 
XU81 n81 n12 VDD VSS INV_X1 
XU80 n12 data_in[34] n19 n86 VDD VSS AOI21_X1 
XU79 n76 n1 VDD VSS INV_X1 
XU78 n1 data_in[50] n10 n92 VDD VSS AOI21_X1 
XU77 data_in[39] n17 VDD VSS INV_X1 
XU75 n77 data_in[38] n17 n87 VDD VSS AOI21_X1 
XU74 data_in[55] n8 VDD VSS INV_X1 
XU73 n72 data_in[54] n8 n93 VDD VSS AOI21_X1 
XU72 n66 n21 VDD VSS INV_X1 
XU71 n23 data_in[15] n21 data_in[19] n65 VDD VSS OAI22_X1 
XU70 n75 n11 n76 n10 n74 VDD VSS AOI22_X1 
XU69 n74 data_in[55] n72 data_in[59] n73 n71 VDD VSS OAI221_X1 
XU68 n80 n20 n81 n19 n79 VDD VSS AOI22_X1 
XU67 n79 data_in[39] n77 data_in[43] n78 n70 VDD VSS OAI221_X1 
XU66 n68 data_in[11] n36 n111 VDD VSS OAI21_X1 
XU65 n102 n103 n104 n105 n101 VDD VSS NAND4_X1 
XU64 n109 n110 n111 n112 n100 VDD VSS NAND4_X1 
XU63 n48 n100 n101 n22 n82 VDD VSS AOI22_X1 
XU62 n113 data_in[4] n33 n69 VDD VSS NOR3_X1 
XU61 n90 data_in[36] n14 n81 VDD VSS NOR3_X1 
XU60 n96 data_in[52] n5 n76 VDD VSS NOR3_X1 
XU59 n54 data_in[8] n34 n67 VDD VSS NOR3_X1 
XU58 n53 data_in[24] n25 n63 VDD VSS NOR3_X1 
XU57 n107 data_in[20] n24 n66 VDD VSS NOR3_X1 
XU56 data_in[16] n30 n24 n106 VDD VSS NOR3_X1 
XU55 data_in[48] n9 n5 n75 VDD VSS NOR3_X1 
XU54 data_in[58] data_in[57] data_in[60] data_in[59] n95 VDD VSS NOR4_X1 
XU53 data_in[42] data_in[41] data_in[44] data_in[43] n89 VDD VSS NOR4_X1 
XU52 data_in[32] n18 n14 n80 VDD VSS NOR3_X1 
XU51 data_in[29] data_in[31] data_in[30] n97 VDD VSS NOR3_X1 
XU50 n80 n55 n97 n47 VDD VSS NAND3_X1 
XU49 data_in[26] data_in[25] data_in[28] data_in[27] n108 VDD VSS NOR4_X1 
XU48 data_in[11] data_in[10] data_in[9] data_in[12] n114 VDD VSS NOR4_X1 
XU47 data_in[34] data_in[33] data_in[36] data_in[35] n90 VDD VSS NOR4_X1 
XU46 data_in[50] data_in[49] data_in[52] data_in[51] n96 VDD VSS NOR4_X1 
XU45 data_in[18] data_in[17] data_in[20] data_in[19] n107 VDD VSS NOR4_X1 
XU43 data_in[21] n25 n116 VDD VSS OR2_X1 
XU42 data_in[23] data_in[24] data_in[22] n116 n53 VDD VSS NOR4_X1 
XU41 data_in[5] n34 n115 VDD VSS OR2_X1 
XU40 data_in[7] data_in[8] data_in[6] n115 n54 VDD VSS NOR4_X1 
XU39 data_in[53] n6 n98 VDD VSS OR2_X1 
XU38 n113 n39 VDD VSS INV_X1 
XU37 n75 n4 VDD VSS INV_X1 
XU36 n106 n23 VDD VSS INV_X1 
XU35 n90 n18 VDD VSS INV_X1 
XU34 n96 n9 VDD VSS INV_X1 
XU33 n107 n30 VDD VSS INV_X1 
XU32 n95 n6 VDD VSS INV_X1 
XU31 n89 n15 VDD VSS INV_X1 
XU30 n108 n25 VDD VSS INV_X1 
XU29 n114 n34 VDD VSS INV_X1 
XU28 n130 data_out[5] VDD VSS INV_X1 
XU27 n53 n25 n30 n24 n52 VDD VSS OAI22_X1 
XU26 n45 n6 n9 n5 n57 VDD VSS OAI22_X1 
XU25 n58 n14 VDD VSS INV_X1 
XU24 n54 n33 VDD VSS INV_X1 
XU23 n53 n24 VDD VSS INV_X1 
XU122 data_in[10] n36 VDD VSS INV_X1 
XU121 data_in[7] n37 VDD VSS INV_X1 
XU120 data_in[11] n35 VDD VSS INV_X1 
XU119 data_in[3] n40 VDD VSS INV_X1 
XU118 data_in[31] n20 VDD VSS INV_X1 
XU1 n131 n3 VDD VSS INV_X1 
XU123 n3 data_out[3] VDD VSS INV_X32 
XU124 n134 n118 VDD VSS INV_X1 
XU125 n118 n119 VDD VSS INV_X32 
XU126 n119 n120 VDD VSS INV_X1 
XU127 n120 data_out[2] VDD VSS INV_X32 
XU128 n133 n122 VDD VSS INV_X1 
XU129 n122 n123 VDD VSS INV_X32 
XU130 n123 n124 VDD VSS INV_X1 
XU131 n124 data_out[1] VDD VSS INV_X32 
XU132 n127 n126 VDD VSS CLKBUF_X1 
XU133 n132 n127 VDD VSS INV_X1 
XU134 n126 data_out[0] VDD VSS INV_X32 
XU135 n47 n129 VDD VSS INV_X32 
XU136 n129 n130 VDD VSS INV_X1 
.ENDS

.SUBCKT gng_coef c2[16] c2[15] c2[14] c2[13] c2[12] c2[11] c2[10] c2[9] c2[8] c2[7] 
+ c2[6] c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] clk VDD VSS c1[17] c1[16] c1[15] c1[14] 
+ c1[13] c1[12] c1[11] c1[10] c1[9] c1[8] c1[7] c1[6] c1[5] c1[4] c1[3] c1[2] c1[1] 
+ c1[0] c0[17] c0[16] c0[15] c0[14] c0[13] c0[12] c0[11] c0[10] c0[9] c0[8] c0[7] 
+ c0[6] c0[5] c0[4] c0[3] c0[2] c0[1] c0[0] addr[7] addr[6] addr[5] addr[4] addr[3] 
+ addr[2] addr[1] addr[0] IN0 IN1 IN2 IN3 IN4 IN5 clk_cts_0 clk_cts_1 
XU1834 n488 n492 n1547 VDD VSS XOR2_X1 
XU1832 n537 n1545 VDD VSS INV_X1 
XU1831 n548 n1544 VDD VSS INV_X1 
XU1830 n539 n1543 VDD VSS INV_X1 
XU1829 n601 n1542 VDD VSS INV_X1 
XU1828 n627 n1541 VDD VSS INV_X1 
XU1827 n6 n1540 VDD VSS INV_X1 
XU1826 n525 n1539 VDD VSS INV_X1 
XU1825 n536 n1538 VDD VSS INV_X1 
XU1824 n1 n1537 VDD VSS INV_X1 
XU1637 addr[0] n515 VDD VSS BUF_X2 
XU1635 addr[0] n513 VDD VSS BUF_X1 
XU1631 addr[0] n509 VDD VSS BUF_X2 
XU1629 addr[1] n507 VDD VSS BUF_X2 
XU1625 addr[1] n503 VDD VSS BUF_X2 
XU1624 addr[1] n502 VDD VSS BUF_X2 
XU1622 addr[1] n500 VDD VSS BUF_X2 
XU1621 addr[1] n499 VDD VSS BUF_X2 
XU1619 addr[1] n497 VDD VSS BUF_X1 
XU1617 addr[1] n495 VDD VSS BUF_X1 
XU1615 IN0 n492 VDD VSS CLKBUF_X2 
XU1597 IN1 n487 VDD VSS BUF_X2 
XU1595 IN1 n484 VDD VSS BUF_X2 
XU1591 IN1 n480 VDD VSS BUF_X2 
XU822 IN2 n477 VDD VSS BUF_X2 
XU707 IN2 n475 VDD VSS BUF_X2 
XU568 IN2 n473 VDD VSS BUF_X2 
XU534 IN2 n471 VDD VSS BUF_X1 
XU521 IN2 n468 VDD VSS BUF_X1 
XU504 IN2 n466 VDD VSS BUF_X2 
XU497 IN2 n464 VDD VSS BUF_X2 
XU491 IN2 n462 VDD VSS BUF_X2 
XU486 IN2 n460 VDD VSS BUF_X2 
XU484 IN2 n458 VDD VSS BUF_X2 
XU481 IN3 n455 VDD VSS BUF_X1 
XU259 IN3 n454 VDD VSS BUF_X2 
XU201 IN3 n453 VDD VSS BUF_X2 
XU147 IN3 n452 VDD VSS BUF_X2 
XU49 IN3 n448 VDD VSS BUF_X2 
XU46 IN4 n445 VDD VSS BUF_X2 
XU28 IN4 n443 VDD VSS BUF_X2 
XU17 IN4 n442 VDD VSS BUF_X2 
XU12 IN4 n439 VDD VSS BUF_X2 
XU10 IN5 n435 VDD VSS BUF_X2 
XU2 n433 n434 VDD VSS INV_X1 
XU1 IN5 n433 VDD VSS BUF_X2 
XU66 n444 n14 n66 VDD VSS XOR2_X1 
XU65 n480 n458 n65 VDD VSS XOR2_X1 
XU64 n493 n1524 n64 VDD VSS XOR2_X1 
XU63 n493 n1536 n63 VDD VSS XOR2_X1 
XU62 n451 n1531 n62 VDD VSS XOR2_X1 
XU61 n488 n497 n61 VDD VSS XOR2_X1 
XU60 n468 n448 n60 VDD VSS XOR2_X1 
XU59 n1531 n1524 addr[5] n59 VDD VSS MUX2_X1 
XU57 n1531 addr[0] n448 n56 VDD VSS MUX2_X1 
XU54 n2 n1 addr[5] n53 VDD VSS MUX2_X1 
XU52 n1531 n1540 addr[5] n51 VDD VSS MUX2_X1 
XU51 n2 addr[0] addr[5] n50 VDD VSS MUX2_X1 
XU50 n6 n2 addr[5] n49 VDD VSS MUX2_X1 
XU48 n9 n1537 addr[5] n47 VDD VSS MUX2_X1 
XU45 n1540 n1524 addr[5] n44 VDD VSS MUX2_X1 
XU43 n1540 n501 n448 n42 VDD VSS MUX2_X1 
XU42 n1 n5 addr[5] n41 VDD VSS MUX2_X1 
XU41 n512 n1540 addr[5] n40 VDD VSS MUX2_X1 
XU40 addr[0] n1524 addr[5] n39 VDD VSS MUX2_X1 
XU38 n1540 n512 addr[5] n37 VDD VSS MUX2_X1 
XU36 n451 addr[1] n35 VDD VSS XOR2_X1 
XU35 n1531 n501 addr[5] n34 VDD VSS MUX2_X1 
XU34 addr[1] n1524 addr[5] n33 VDD VSS MUX2_X1 
XU33 n1524 n501 addr[5] n32 VDD VSS MUX2_X1 
XU32 n1531 addr[1] addr[5] n31 VDD VSS MUX2_X1 
XU31 n9 addr[0] addr[5] n30 VDD VSS MUX2_X1 
XU29 n2 addr[5] n28 VDD VSS XOR2_X1 
XU27 addr[0] n497 n448 n26 VDD VSS MUX2_X1 
XU26 n1537 n512 n448 n25 VDD VSS MUX2_X1 
XU25 n1537 addr[0] n448 n24 VDD VSS MUX2_X1 
XU24 n512 n2 n448 n23 VDD VSS MUX2_X1 
XU23 addr[0] n2 n448 n22 VDD VSS MUX2_X1 
XU21 n1527 addr[1] addr[5] n20 VDD VSS MUX2_X1 
XU19 n5 n501 n448 n18 VDD VSS MUX2_X1 
XU16 n501 addr[0] n9 VDD VSS XOR2_X1 
XU15 n1537 n1527 n448 n17 VDD VSS MUX2_X1 
Xc1_reg_0_ d[17] n63_G2B1I9 n2037 SYNOPSYS_UNCONNECTED_272 VDD VSS DFF_X1 
Xc1_reg_1_ d[18] n63_G2B1I9 n2038 SYNOPSYS_UNCONNECTED_271 VDD VSS DFF_X1 
Xc1_reg_2_ d[19] n63_G2B1I9 n2039 SYNOPSYS_UNCONNECTED_270 VDD VSS DFF_X1 
Xc1_reg_3_ d[20] n63_G2B1I9 n2040 SYNOPSYS_UNCONNECTED_269 VDD VSS DFF_X1 
Xc1_reg_4_ d[21] n63_G2B1I9 n2041 SYNOPSYS_UNCONNECTED_268 VDD VSS DFF_X1 
Xc1_reg_5_ d[22] n63_G2B1I7 n2042 SYNOPSYS_UNCONNECTED_267 VDD VSS DFF_X1 
Xc1_reg_6_ d[23] n63_G2B1I7 n2027 SYNOPSYS_UNCONNECTED_266 VDD VSS DFF_X1 
Xc1_reg_7_ d[24] n63_G2B1I7 n2028 SYNOPSYS_UNCONNECTED_265 VDD VSS DFF_X1 
Xc1_reg_8_ d[25] n63_G2B1I7 n2029 SYNOPSYS_UNCONNECTED_264 VDD VSS DFF_X1 
Xc1_reg_9_ d[26] n63_G2B1I7 n2030 SYNOPSYS_UNCONNECTED_263 VDD VSS DFF_X1 
Xc1_reg_10_ d[27] n63_G2B1I7 n2031 SYNOPSYS_UNCONNECTED_262 VDD VSS DFF_X1 
Xc1_reg_11_ d[28] n63_G2B1I7 n2032 SYNOPSYS_UNCONNECTED_261 VDD VSS DFF_X1 
Xc1_reg_12_ n457 clk_cts_1 n2033 SYNOPSYS_UNCONNECTED_260 VDD VSS DFF_X1 
Xc1_reg_13_ d[30] clk_cts_1 n2034 SYNOPSYS_UNCONNECTED_259 VDD VSS DFF_X1 
Xc1_reg_14_ n1548 clk_cts_0 n2019 SYNOPSYS_UNCONNECTED_258 VDD VSS DFF_X1 
Xc1_reg_15_ n514 clk_cts_0 n2020 SYNOPSYS_UNCONNECTED_257 VDD VSS DFF_X1 
Xc1_reg_16_ n2061 clk_cts_0 n2021 SYNOPSYS_UNCONNECTED_256 VDD VSS DFF_X1 
Xc0_reg_0_ d[35] n63_G2B1I6 n2051 SYNOPSYS_UNCONNECTED_255 VDD VSS DFF_X1 
Xc0_reg_1_ d[36] n63_G2B1I6 n2052 SYNOPSYS_UNCONNECTED_254 VDD VSS DFF_X1 
Xc0_reg_2_ d[37] n63_G2B1I6 n2053 SYNOPSYS_UNCONNECTED_253 VDD VSS DFF_X1 
Xc0_reg_3_ d[38] n63_G2B1I6 n2054 SYNOPSYS_UNCONNECTED_252 VDD VSS DFF_X1 
Xc0_reg_4_ d[39] n63_G2B1I5 n2055 SYNOPSYS_UNCONNECTED_251 VDD VSS DFF_X1 
Xc0_reg_5_ d[40] n63_G2B1I5 n2056 SYNOPSYS_UNCONNECTED_250 VDD VSS DFF_X1 
Xc0_reg_6_ d[41] n63_G2B1I5 n2057 SYNOPSYS_UNCONNECTED_249 VDD VSS DFF_X1 
Xc0_reg_7_ d[42] n63_G2B1I6 n2058 SYNOPSYS_UNCONNECTED_248 VDD VSS DFF_X1 
Xc0_reg_8_ d[43] n63_G2B1I5 n2043 SYNOPSYS_UNCONNECTED_247 VDD VSS DFF_X1 
Xc0_reg_9_ n506 clk_cts_1 n2044 SYNOPSYS_UNCONNECTED_246 VDD VSS DFF_X1 
Xc0_reg_10_ n504 clk_cts_0 n2045 SYNOPSYS_UNCONNECTED_245 VDD VSS DFF_X1 
Xc0_reg_11_ n498 n63_G2B1I9 n2046 SYNOPSYS_UNCONNECTED_244 VDD VSS DFF_X1 
Xc0_reg_12_ n496 n63_G2B1I9 n2047 SYNOPSYS_UNCONNECTED_243 VDD VSS DFF_X1 
Xc0_reg_13_ n494 n63_G2B1I9 n2048 SYNOPSYS_UNCONNECTED_242 VDD VSS DFF_X1 
Xc0_reg_14_ n490 n63_G2B1I6 n2049 SYNOPSYS_UNCONNECTED_241 VDD VSS DFF_X1 
Xc0_reg_15_ n2060 n63_G2B1I1 n2050 SYNOPSYS_UNCONNECTED_240 VDD VSS DFF_X1 
Xc0_reg_16_ N4680 n63_G2B1I6 n2035 SYNOPSYS_UNCONNECTED_239 VDD VSS DFF_X1 
Xc0_reg_17_ N4640 n63_G2B1I1 n2036 SYNOPSYS_UNCONNECTED_238 VDD VSS DFF_X1 
Xc2_reg_0_ d[0] n63_G2B1I4 n2023 SYNOPSYS_UNCONNECTED_237 VDD VSS DFF_X1 
Xc2_reg_1_ d[1] clk_cts_0 n2024 SYNOPSYS_UNCONNECTED_236 VDD VSS DFF_X1 
Xc2_reg_2_ d[2] n63_G2B1I1 n2025 SYNOPSYS_UNCONNECTED_235 VDD VSS DFF_X1 
Xc2_reg_3_ d[3] n63_G2B1I9 n2026 SYNOPSYS_UNCONNECTED_234 VDD VSS DFF_X1 
Xc2_reg_4_ d[4] n63_G2B1I3 n2011 SYNOPSYS_UNCONNECTED_233 VDD VSS DFF_X1 
Xc2_reg_5_ n478 n63_G2B1I3 n2012 SYNOPSYS_UNCONNECTED_232 VDD VSS DFF_X1 
Xc2_reg_6_ n474 n63_G2B1I3 n2013 SYNOPSYS_UNCONNECTED_231 VDD VSS DFF_X1 
Xc2_reg_7_ d[7] n63_G2B1I1 n2014 SYNOPSYS_UNCONNECTED_230 VDD VSS DFF_X1 
Xc2_reg_8_ n470 n63_G2B1I3 n2015 SYNOPSYS_UNCONNECTED_229 VDD VSS DFF_X1 
Xc2_reg_9_ n467 n63_G2B1I3 n2016 SYNOPSYS_UNCONNECTED_228 VDD VSS DFF_X1 
Xc2_reg_10_ d[10] n63_G2B1I4 n2017 SYNOPSYS_UNCONNECTED_227 VDD VSS DFF_X1 
Xc2_reg_11_ d[11] n63_G2B1I4 n2018 SYNOPSYS_UNCONNECTED_226 VDD VSS DFF_X1 
Xc2_reg_12_ d[12] n63_G2B1I4 n2006 SYNOPSYS_UNCONNECTED_225 VDD VSS DFF_X1 
Xc2_reg_13_ d[13] n63_G2B1I4 n2007 SYNOPSYS_UNCONNECTED_224 VDD VSS DFF_X1 
Xc2_reg_14_ d[14] n63_G2B1I4 n2008 SYNOPSYS_UNCONNECTED_223 VDD VSS DFF_X1 
Xc2_reg_15_ n459 n63_G2B1I4 n2009 SYNOPSYS_UNCONNECTED_222 VDD VSS DFF_X1 
Xc2_reg_16_ N19520 n63_G2B1I4 n2010 SYNOPSYS_UNCONNECTED_221 VDD VSS DFF_X1 
XU162 n160 n151 addr[7] n161 VDD VSS MUX2_X1 
XU161 n159 n155 addr[4] n160 VDD VSS MUX2_X1 
XU160 n158 n156 addr[3] n159 VDD VSS MUX2_X1 
XU159 n157 n1630 addr[2] n158 VDD VSS MUX2_X1 
XU158 n1 addr[1] addr[5] n157 VDD VSS MUX2_X1 
XU157 n1631 n1632 addr[2] n156 VDD VSS MUX2_X1 
XU156 n154 n152 addr[3] n155 VDD VSS MUX2_X1 
XU155 n153 n62 addr[2] n154 VDD VSS MUX2_X1 
XU154 n2 addr[1] addr[5] n153 VDD VSS MUX2_X1 
XU153 n1648 n1628 addr[2] n152 VDD VSS MUX2_X1 
XU152 n150 n147 addr[4] n151 VDD VSS MUX2_X1 
XU151 n149 n148 n484 n150 VDD VSS MUX2_X1 
XU150 n11 n1597 addr[2] n149 VDD VSS MUX2_X1 
XU149 n32 n5 addr[2] n148 VDD VSS MUX2_X1 
XU148 n146 n145 n484 n147 VDD VSS MUX2_X1 
XU146 addr[1] n1596 IN0 n145 VDD VSS MUX2_X1 
XU145 n143 n138 addr[7] n144 VDD VSS MUX2_X1 
XU144 n142 n140 n458 n143 VDD VSS MUX2_X1 
XU143 n141 n64 n484 n142 VDD VSS MUX2_X1 
XU142 n1633 n1634 IN0 n141 VDD VSS MUX2_X1 
XU141 n139 n63 n484 n140 VDD VSS MUX2_X1 
XU140 n5 n1596 IN0 n139 VDD VSS MUX2_X1 
XU139 n137 n135 n458 n138 VDD VSS MUX2_X1 
XU138 n449 n136 n429 n137 VDD VSS MUX2_X1 
XU137 n12 n411 n480 n136 VDD VSS MUX2_X1 
XU136 n134 n1598 n484 n135 VDD VSS MUX2_X1 
XU135 n1655 n430 IN0 n134 VDD VSS MUX2_X1 
XU134 n133 n116 addr[6] d[45] VDD VSS MUX2_X1 
XU133 n132 n123 addr[7] n133 VDD VSS MUX2_X1 
XU132 n131 n126 addr[4] n132 VDD VSS MUX2_X1 
XU131 n128 n129 addr[2] n131 VDD VSS MUX2_X1 
XU129 n1624 n127 addr[3] n128 VDD VSS MUX2_X1 
XU128 addr[1] n9 addr[5] n127 VDD VSS MUX2_X1 
XU127 n125 n124 IN0 n126 VDD VSS MUX2_X1 
XU126 n1645 n1651 n487 n125 VDD VSS MUX2_X1 
XU125 addr[0] n22 n487 n124 VDD VSS MUX2_X1 
XU124 n122 n119 addr[4] n123 VDD VSS MUX2_X1 
XU123 n121 n120 addr[2] n122 VDD VSS MUX2_X1 
XU122 n1625 n1626 addr[3] n121 VDD VSS MUX2_X1 
XU121 n33 n8 addr[3] n120 VDD VSS MUX2_X1 
XU120 n61 n118 IN0 n119 VDD VSS MUX2_X1 
XU119 n9 n117 n484 n118 VDD VSS MUX2_X1 
XU118 n5 n6 n448 n117 VDD VSS MUX2_X1 
XU117 n115 n108 addr[7] n116 VDD VSS MUX2_X1 
XU116 n114 n111 addr[4] n115 VDD VSS MUX2_X1 
XU115 n113 n112 addr[2] n114 VDD VSS MUX2_X1 
XU114 n1628 n27 addr[3] n113 VDD VSS MUX2_X1 
XU113 n1627 n1531 addr[3] n112 VDD VSS MUX2_X1 
XU112 n110 n109 addr[2] n111 VDD VSS MUX2_X1 
XU111 n1531 n1595 addr[3] n110 VDD VSS MUX2_X1 
XU110 n34 n33 addr[3] n109 VDD VSS MUX2_X1 
XU109 n107 n103 addr[4] n108 VDD VSS MUX2_X1 
XU108 n106 n104 addr[2] n107 VDD VSS MUX2_X1 
XU107 n105 n8 addr[3] n106 VDD VSS MUX2_X1 
XU105 n33 n32 addr[3] n104 VDD VSS MUX2_X1 
XU104 n102 n101 addr[2] n103 VDD VSS MUX2_X1 
XU103 n1654 n1596 n484 n102 VDD VSS MUX2_X1 
XU102 n1629 n1597 n484 n101 VDD VSS MUX2_X1 
XU101 n100 n83 n445 d[44] VDD VSS MUX2_X1 
XU100 n99 n91 n433 n100 VDD VSS MUX2_X1 
XU99 n98 n94 IN0 n99 VDD VSS MUX2_X1 
XU98 n97 n95 n487 n98 VDD VSS MUX2_X1 
XU97 n1609 n96 n460 n97 VDD VSS MUX2_X1 
XU96 n497 n1531 n448 n96 VDD VSS MUX2_X1 
XU95 n1653 n3 n460 n95 VDD VSS MUX2_X1 
XU94 n93 n92 n487 n94 VDD VSS MUX2_X1 
XU93 n1614 n1613 n460 n93 VDD VSS MUX2_X1 
XU92 n1616 n1617 n460 n92 VDD VSS MUX2_X1 
XU91 n90 n86 IN0 n91 VDD VSS MUX2_X1 
XU90 n89 n88 n487 n90 VDD VSS MUX2_X1 
XU89 n22 n23 n460 n89 VDD VSS MUX2_X1 
XU88 n87 n2 n60 n88 VDD VSS MUX2_X1 
XU87 n1527 n512 n468 n87 VDD VSS MUX2_X1 
XU86 n85 n84 n487 n86 VDD VSS MUX2_X1 
XU85 n1618 addr[0] n460 n85 VDD VSS MUX2_X1 
XU84 n1619 n1652 n460 n84 VDD VSS MUX2_X1 
XU83 n82 n75 n433 n83 VDD VSS MUX2_X1 
XU82 n81 n78 IN0 n82 VDD VSS MUX2_X1 
XU81 n80 n79 n487 n81 VDD VSS MUX2_X1 
XU80 n1620 n1621 n460 n80 VDD VSS MUX2_X1 
XU79 n24 n512 n460 n79 VDD VSS MUX2_X1 
XU78 n77 n76 n487 n78 VDD VSS MUX2_X1 
XU77 n1622 n1620 n460 n77 VDD VSS MUX2_X1 
XU76 addr[0] n1618 n460 n76 VDD VSS MUX2_X1 
XU75 n74 n71 IN0 n75 VDD VSS MUX2_X1 
XU74 n73 n72 n487 n74 VDD VSS MUX2_X1 
XU73 n1652 n1607 n460 n73 VDD VSS MUX2_X1 
XU72 n1651 n1602 n468 n72 VDD VSS MUX2_X1 
XU71 n1604 n70 n487 n71 VDD VSS MUX2_X1 
XU70 n1645 n1594 n460 n70 VDD VSS MUX2_X1 
XU69 n449 n1 n69 VDD VSS XOR2_X1 
XU68 n448 n433 n68 VDD VSS XOR2_X1 
XU67 n480 n433 n67 VDD VSS XOR2_X1 
XU273 n27 n271 n433 n272 VDD VSS MUX2_X1 
XU272 n501 n1537 n448 n271 VDD VSS MUX2_X1 
XU271 n269 n1524 n68 n270 VDD VSS MUX2_X1 
XU270 n5 n1537 n433 n269 VDD VSS MUX2_X1 
XU269 n267 n266 n487 n268 VDD VSS MUX2_X1 
XU267 n1658 n26 addr[7] n266 VDD VSS MUX2_X1 
XU266 n264 n260 addr[2] n265 VDD VSS MUX2_X1 
XU265 n263 n262 n487 n264 VDD VSS MUX2_X1 
XU264 n47 n1 addr[7] n263 VDD VSS MUX2_X1 
XU263 n58 n261 addr[7] n262 VDD VSS MUX2_X1 
XU260 n258 n259 n487 n260 VDD VSS MUX2_X1 
XU258 n1656 n1657 addr[7] n258 VDD VSS MUX2_X1 
XU257 n256 n250 n460 n257 VDD VSS MUX2_X1 
XU256 n255 n253 n492 n256 VDD VSS MUX2_X1 
XU255 n254 n1655 n67 n255 VDD VSS MUX2_X1 
XU254 n43 n1640 n484 n254 VDD VSS MUX2_X1 
XU253 n252 n251 n487 n253 VDD VSS MUX2_X1 
XU251 n1615 n1536 n433 n251 VDD VSS MUX2_X1 
XU250 n249 n245 IN0 n250 VDD VSS MUX2_X1 
XU249 n247 n246 n484 n249 VDD VSS MUX2_X1 
XU247 n1650 n1597 addr[7] n246 VDD VSS MUX2_X1 
XU246 n244 n242 n484 n245 VDD VSS MUX2_X1 
XU245 n243 n1605 addr[7] n244 VDD VSS MUX2_X1 
XU244 n501 n1524 n455 n243 VDD VSS MUX2_X1 
XU243 n1606 n1591 addr[7] n242 VDD VSS MUX2_X1 
XU242 n241 n225 addr[6] d[4] VDD VSS MUX2_X1 
XU241 n240 n232 addr[7] n241 VDD VSS MUX2_X1 
XU240 n239 n234 addr[4] n240 VDD VSS MUX2_X1 
XU239 n238 n237 addr[2] n239 VDD VSS MUX2_X1 
XU238 n1631 n1637 addr[3] n238 VDD VSS MUX2_X1 
XU237 n236 n235 addr[3] n237 VDD VSS MUX2_X1 
XU236 n2 n6 addr[5] n236 VDD VSS MUX2_X1 
XU235 n1527 n1524 addr[5] n235 VDD VSS MUX2_X1 
XU234 n233 n1597 addr[2] n234 VDD VSS MUX2_X1 
XU233 n1611 n512 n487 n233 VDD VSS MUX2_X1 
XU232 n231 n228 addr[4] n232 VDD VSS MUX2_X1 
XU231 n230 n229 addr[2] n231 VDD VSS MUX2_X1 
XU230 n37 n15 addr[3] n230 VDD VSS MUX2_X1 
XU229 n26 n39 addr[3] n229 VDD VSS MUX2_X1 
XU228 n227 n226 addr[2] n228 VDD VSS MUX2_X1 
XU227 n411 n1638 n487 n227 VDD VSS MUX2_X1 
XU226 n30 n1639 addr[3] n226 VDD VSS MUX2_X1 
XU225 n224 n216 addr[7] n225 VDD VSS MUX2_X1 
XU224 n222 n219 addr[4] n224 VDD VSS MUX2_X1 
XU222 n221 n1611 addr[2] n220 VDD VSS MUX2_X1 
XU221 n218 n217 addr[2] n219 VDD VSS MUX2_X1 
XU220 n7 n1640 addr[3] n218 VDD VSS MUX2_X1 
XU219 n6 n1599 n484 n217 VDD VSS MUX2_X1 
XU218 n215 n212 addr[4] n216 VDD VSS MUX2_X1 
XU217 n214 n213 addr[2] n215 VDD VSS MUX2_X1 
XU216 n427 n1591 n484 n214 VDD VSS MUX2_X1 
XU215 n105 n1594 n484 n213 VDD VSS MUX2_X1 
XU214 n211 n210 n492 n212 VDD VSS MUX2_X1 
XU212 n1605 n449 n484 n210 VDD VSS MUX2_X1 
XU211 n209 n196 addr[7] d[48] VDD VSS MUX2_X1 
XU210 n208 n202 n458 n209 VDD VSS MUX2_X1 
XU209 n206 n207 IN0 n208 VDD VSS MUX2_X1 
XU207 n205 n203 n445 n206 VDD VSS MUX2_X1 
XU204 n199 n200 IN0 n202 VDD VSS MUX2_X1 
XU202 n197 n198 n445 n199 VDD VSS MUX2_X1 
XU200 n12 n427 n480 n197 VDD VSS MUX2_X1 
XU199 n195 n191 n458 n196 VDD VSS MUX2_X1 
XU198 n66 n194 IN0 n195 VDD VSS MUX2_X1 
XU197 n193 n192 n445 n194 VDD VSS MUX2_X1 
XU195 n12 n455 n480 n192 VDD VSS MUX2_X1 
XU194 n190 n187 IN0 n191 VDD VSS MUX2_X1 
XU193 n189 n188 n445 n190 VDD VSS MUX2_X1 
XU190 n14 n186 n445 n187 VDD VSS MUX2_X1 
XU189 n1636 n1536 n484 n186 VDD VSS MUX2_X1 
XU188 n185 n171 n445 d[47] VDD VSS MUX2_X1 
XU187 n184 n177 addr[7] n185 VDD VSS MUX2_X1 
XU186 n183 n180 addr[4] n184 VDD VSS MUX2_X1 
XU185 n182 n181 n484 n183 VDD VSS MUX2_X1 
XU184 n31 n33 addr[2] n182 VDD VSS MUX2_X1 
XU183 n13 n1536 IN0 n181 VDD VSS MUX2_X1 
XU182 n179 n178 n484 n180 VDD VSS MUX2_X1 
XU181 n1595 n1635 addr[2] n179 VDD VSS MUX2_X1 
XU180 n1591 n1656 addr[2] n178 VDD VSS MUX2_X1 
XU179 n176 n173 n458 n177 VDD VSS MUX2_X1 
XU178 n175 n174 n480 n176 VDD VSS MUX2_X1 
XU177 n449 n12 IN0 n175 VDD VSS MUX2_X1 
XU176 n455 n411 IN0 n174 VDD VSS MUX2_X1 
XU175 n449 n172 n484 n173 VDD VSS MUX2_X1 
XU174 n1595 n455 IN0 n172 VDD VSS MUX2_X1 
XU173 n170 n165 addr[7] n171 VDD VSS MUX2_X1 
XU172 n169 n167 n458 n170 VDD VSS MUX2_X1 
XU171 n168 n45 n480 n169 VDD VSS MUX2_X1 
XU169 n1851 n166 n480 n167 VDD VSS MUX2_X1 
XU167 n1598 n164 n65 n165 VDD VSS MUX2_X1 
XU166 n163 n162 n458 n164 VDD VSS MUX2_X1 
XU165 n1634 n455 n492 n163 VDD VSS MUX2_X1 
XU164 n38 n19 n492 n162 VDD VSS MUX2_X1 
XU163 n161 n144 addr[6] d[46] VDD VSS MUX2_X1 
XU376 n374 n366 n460 n375 VDD VSS MUX2_X1 
XU375 n373 n369 addr[2] n374 VDD VSS MUX2_X1 
XU374 n372 n370 n487 n373 VDD VSS MUX2_X1 
XU373 n16 n371 addr[7] n372 VDD VSS MUX2_X1 
XU372 addr[0] n1540 addr[5] n371 VDD VSS MUX2_X1 
XU371 addr[1] n1658 addr[7] n370 VDD VSS MUX2_X1 
XU370 n368 n367 n487 n369 VDD VSS MUX2_X1 
XU369 n9 n46 addr[7] n368 VDD VSS MUX2_X1 
XU368 n1617 n19 addr[7] n367 VDD VSS MUX2_X1 
XU367 n365 n361 addr[2] n366 VDD VSS MUX2_X1 
XU366 n364 n362 n487 n365 VDD VSS MUX2_X1 
XU365 n363 n12 addr[7] n364 VDD VSS MUX2_X1 
XU364 n6 n1 n448 n363 VDD VSS MUX2_X1 
XU363 n3 n1622 addr[7] n362 VDD VSS MUX2_X1 
XU362 n360 n359 n487 n361 VDD VSS MUX2_X1 
XU361 n41 n20 addr[7] n360 VDD VSS MUX2_X1 
XU360 n36 n358 addr[7] n359 VDD VSS MUX2_X1 
XU358 n356 n348 n460 n357 VDD VSS MUX2_X1 
XU357 n355 n352 IN0 n356 VDD VSS MUX2_X1 
XU356 n353 n354 n487 n355 VDD VSS MUX2_X1 
XU354 n1638 n1607 addr[7] n353 VDD VSS MUX2_X1 
XU353 n350 n351 n487 n352 VDD VSS MUX2_X1 
XU351 n52 n349 addr[7] n350 VDD VSS MUX2_X1 
XU350 n5 n9 n448 n349 VDD VSS MUX2_X1 
XU349 n345 n346 IN0 n348 VDD VSS MUX2_X1 
XU347 n344 n343 n484 n345 VDD VSS MUX2_X1 
XU346 n1605 n1599 addr[7] n344 VDD VSS MUX2_X1 
XU345 n56 n342 addr[7] n343 VDD VSS MUX2_X1 
XU343 n430 n69 n480 n341 VDD VSS MUX2_X1 
XU342 n340 n324 addr[6] d[7] VDD VSS MUX2_X1 
XU341 n339 n332 addr[7] n340 VDD VSS MUX2_X1 
XU340 n338 n335 addr[4] n339 VDD VSS MUX2_X1 
XU339 n337 n336 addr[2] n338 VDD VSS MUX2_X1 
XU338 n1603 n31 n484 n337 VDD VSS MUX2_X1 
XU337 n1599 n5 n484 n336 VDD VSS MUX2_X1 
XU336 n334 n333 addr[2] n335 VDD VSS MUX2_X1 
XU335 n56 n1608 n484 n334 VDD VSS MUX2_X1 
XU334 n1634 n1625 n484 n333 VDD VSS MUX2_X1 
XU333 n331 n327 addr[4] n332 VDD VSS MUX2_X1 
XU332 n330 n329 addr[2] n331 VDD VSS MUX2_X1 
XU331 n1625 n1612 n484 n330 VDD VSS MUX2_X1 
XU330 n328 n7 n484 n329 VDD VSS MUX2_X1 
XU328 n326 n325 addr[2] n327 VDD VSS MUX2_X1 
XU327 n1639 n8 addr[3] n326 VDD VSS MUX2_X1 
XU326 n1653 n451 n484 n325 VDD VSS MUX2_X1 
XU325 n323 n313 addr[7] n324 VDD VSS MUX2_X1 
XU324 n322 n318 addr[4] n323 VDD VSS MUX2_X1 
XU323 n321 n319 addr[2] n322 VDD VSS MUX2_X1 
XU322 n512 n320 n484 n321 VDD VSS MUX2_X1 
XU321 n5 addr[0] addr[5] n320 VDD VSS MUX2_X1 
XU320 n25 n51 n484 n319 VDD VSS MUX2_X1 
XU319 n315 n316 addr[2] n318 VDD VSS MUX2_X1 
XU317 n314 n1595 n484 n315 VDD VSS MUX2_X1 
XU316 n512 n1 addr[5] n314 VDD VSS MUX2_X1 
XU315 n312 n307 addr[4] n313 VDD VSS MUX2_X1 
XU314 n309 n310 addr[2] n312 VDD VSS MUX2_X1 
XU312 n1626 n308 n484 n309 VDD VSS MUX2_X1 
XU311 n1537 n9 addr[5] n308 VDD VSS MUX2_X1 
XU310 n306 n305 addr[2] n307 VDD VSS MUX2_X1 
XU308 n1599 n451 n484 n305 VDD VSS MUX2_X1 
XU307 n304 n289 addr[6] d[6] VDD VSS MUX2_X1 
XU306 n303 n296 addr[7] n304 VDD VSS MUX2_X1 
XU305 n302 n299 n460 n303 VDD VSS MUX2_X1 
XU304 n301 n300 IN0 n302 VDD VSS MUX2_X1 
XU303 n1612 n1661 n487 n301 VDD VSS MUX2_X1 
XU302 n1660 n1641 n487 n300 VDD VSS MUX2_X1 
XU301 n298 n297 IN0 n299 VDD VSS MUX2_X1 
XU299 n1610 n54 n487 n297 VDD VSS MUX2_X1 
XU298 n295 n292 n460 n296 VDD VSS MUX2_X1 
XU297 n294 n293 addr[2] n295 VDD VSS MUX2_X1 
XU296 n50 n35 addr[3] n294 VDD VSS MUX2_X1 
XU295 n1637 n16 addr[3] n293 VDD VSS MUX2_X1 
XU294 n291 n290 addr[2] n292 VDD VSS MUX2_X1 
XU293 n15 n1640 addr[3] n291 VDD VSS MUX2_X1 
XU292 n1660 n53 n487 n290 VDD VSS MUX2_X1 
XU291 n288 n281 addr[7] n289 VDD VSS MUX2_X1 
XU290 n287 n284 n460 n288 VDD VSS MUX2_X1 
XU289 n286 n285 IN0 n287 VDD VSS MUX2_X1 
XU288 n1633 n1641 n487 n286 VDD VSS MUX2_X1 
XU287 n21 n4 n487 n285 VDD VSS MUX2_X1 
XU286 n283 n282 IN0 n284 VDD VSS MUX2_X1 
XU285 n1659 n40 n487 n283 VDD VSS MUX2_X1 
XU284 n1594 n1622 n487 n282 VDD VSS MUX2_X1 
XU283 n280 n277 addr[4] n281 VDD VSS MUX2_X1 
XU282 n279 n278 addr[2] n280 VDD VSS MUX2_X1 
XU281 n1625 n1629 addr[3] n279 VDD VSS MUX2_X1 
XU280 n1647 n1594 addr[3] n278 VDD VSS MUX2_X1 
XU279 n1600 n276 n429 n277 VDD VSS MUX2_X1 
XU278 n1591 n1536 n492 n276 VDD VSS MUX2_X1 
XU277 n275 n257 addr[6] d[5] VDD VSS MUX2_X1 
XU276 n274 n265 n460 n275 VDD VSS MUX2_X1 
XU275 n273 n268 addr[2] n274 VDD VSS MUX2_X1 
XU274 n272 n270 n487 n273 VDD VSS MUX2_X1 
XU619 n533 n1520 n515 n608 VDD VSS MUX2_X1 
XU617 n1522 n492 n509 n606 VDD VSS MUX2_X1 
XU616 n1526 n1522 n515 n605 VDD VSS MUX2_X1 
XU614 n517 n1522 n509 n603 VDD VSS MUX2_X1 
XU613 n488 n492 n515 n602 VDD VSS MUX2_X1 
XU612 n1526 n488 n515 n601 VDD VSS MUX2_X1 
XU610 n488 n528 n509 n599 VDD VSS MUX2_X1 
XU609 n492 n480 n513 n598 VDD VSS MUX2_X1 
XU607 n1318 n492 n515 n596 VDD VSS MUX2_X1 
XU606 n526 n492 n509 n595 VDD VSS MUX2_X1 
XU605 n493 n517 n509 n594 VDD VSS MUX2_X1 
XU602 n1318 n1522 n515 n591 VDD VSS MUX2_X1 
XU601 n517 n515 n590 VDD VSS XOR2_X1 
XU600 n492 n1526 n509 n589 VDD VSS MUX2_X1 
XU599 IN1 n526 n515 n588 VDD VSS MUX2_X1 
XU597 n517 n488 n509 n586 VDD VSS MUX2_X1 
XU596 n1525 n1526 n515 n585 VDD VSS MUX2_X1 
XU595 n1525 n492 n509 n584 VDD VSS MUX2_X1 
XU594 n533 n492 n515 n583 VDD VSS MUX2_X1 
XU590 n488 n513 n579 VDD VSS XOR2_X1 
XU589 n520 IN1 n515 n578 VDD VSS MUX2_X1 
XU588 n520 n526 n509 n577 VDD VSS MUX2_X1 
XU587 n492 n1520 n515 n576 VDD VSS MUX2_X1 
XU586 n517 n492 n515 n575 VDD VSS MUX2_X1 
XU584 n488 n533 n515 n573 VDD VSS MUX2_X1 
XU583 n480 n520 n513 n547 VDD VSS MUX2_X1 
XU582 n1520 n1526 n515 n572 VDD VSS MUX2_X1 
XU581 n1522 IN1 n515 n571 VDD VSS MUX2_X1 
XU580 n492 n528 n515 n570 VDD VSS MUX2_X1 
XU578 n449 n468 n568 VDD VSS XOR2_X1 
XU577 n488 n526 n515 n567 VDD VSS MUX2_X1 
XU576 n1526 n1318 n515 n566 VDD VSS MUX2_X1 
XU575 n533 n526 n509 n565 VDD VSS MUX2_X1 
XU574 n492 n1522 n515 n564 VDD VSS MUX2_X1 
XU573 n1522 n517 n509 n563 VDD VSS MUX2_X1 
XU572 IN1 n492 n515 n562 VDD VSS MUX2_X1 
XU571 n512 n1522 n561 VDD VSS XOR2_X1 
XU569 n528 n517 n509 n559 VDD VSS MUX2_X1 
XU567 n533 IN1 n515 n557 VDD VSS MUX2_X1 
XU566 n528 n520 n509 n556 VDD VSS MUX2_X1 
XU564 n488 n1522 n509 n554 VDD VSS MUX2_X1 
XU563 n1318 n1525 n515 n553 VDD VSS MUX2_X1 
XU557 n1520 n533 n509 n550 VDD VSS MUX2_X1 
XU556 n493 n1318 n509 n549 VDD VSS MUX2_X1 
XU554 n488 n492 n533 VDD VSS XOR2_X1 
XU439 n1614 n1610 n487 n402 VDD VSS MUX2_X1 
XU438 n426 n461 n487 n403 VDD VSS MUX2_X1 
XU436 addr[0] n9 n448 n425 VDD VSS MUX2_X1 
XU435 n406 n13 n480 n347 VDD VSS MUX2_X1 
XU434 addr[0] n1 n448 n424 VDD VSS MUX2_X1 
XU433 n501 n1 n448 n423 VDD VSS MUX2_X1 
XU432 n1540 n1531 addr[5] n422 VDD VSS MUX2_X1 
XU431 n5 n2 addr[5] n421 VDD VSS MUX2_X1 
XU430 addr[1] n2 addr[5] n420 VDD VSS MUX2_X1 
XU429 n41 n43 addr[2] n223 VDD VSS MUX2_X1 
XU428 n1646 n449 n480 n201 VDD VSS MUX2_X1 
XU427 n1540 addr[1] addr[5] n419 VDD VSS MUX2_X1 
XU426 n501 n1540 n448 n418 VDD VSS MUX2_X1 
XU425 n455 n38 IN0 n417 VDD VSS MUX2_X1 
XU424 n501 n6 n448 n416 VDD VSS MUX2_X1 
XU423 n1537 addr[1] addr[5] n415 VDD VSS MUX2_X1 
XU422 n2 n1531 n448 n414 VDD VSS MUX2_X1 
XU421 n512 n9 n448 n413 VDD VSS MUX2_X1 
XU420 n1623 n407 n460 n412 VDD VSS MUX2_X1 
XU407 n9 n1527 addr[5] n221 VDD VSS MUX2_X1 
XU406 n405 n389 addr[6] d[9] VDD VSS MUX2_X1 
XU405 n404 n397 addr[7] n405 VDD VSS MUX2_X1 
XU404 n400 n401 IN0 n404 VDD VSS MUX2_X1 
XU402 n399 n398 n487 n400 VDD VSS MUX2_X1 
XU401 n1 n1644 n460 n399 VDD VSS MUX2_X1 
XU400 n41 n1662 n460 n398 VDD VSS MUX2_X1 
XU399 n396 n392 IN0 n397 VDD VSS MUX2_X1 
XU398 n395 n393 n484 n396 VDD VSS MUX2_X1 
XU397 n1654 n394 addr[4] n395 VDD VSS MUX2_X1 
XU396 n512 n1524 addr[5] n394 VDD VSS MUX2_X1 
XU395 n52 n1657 addr[4] n393 VDD VSS MUX2_X1 
XU394 n391 n390 n487 n392 VDD VSS MUX2_X1 
XU393 n55 n59 n460 n391 VDD VSS MUX2_X1 
XU392 n1662 n1638 n460 n390 VDD VSS MUX2_X1 
XU391 n388 n381 addr[7] n389 VDD VSS MUX2_X1 
XU390 n387 n384 addr[2] n388 VDD VSS MUX2_X1 
XU389 n386 n385 n487 n387 VDD VSS MUX2_X1 
XU388 n57 n1642 n460 n386 VDD VSS MUX2_X1 
XU387 n1536 n1649 n460 n385 VDD VSS MUX2_X1 
XU386 n383 n382 n487 n384 VDD VSS MUX2_X1 
XU385 n1616 n1659 n460 n383 VDD VSS MUX2_X1 
XU384 n49 n1631 n460 n382 VDD VSS MUX2_X1 
XU383 n380 n377 addr[2] n381 VDD VSS MUX2_X1 
XU382 n379 n378 n487 n380 VDD VSS MUX2_X1 
XU380 n1595 n1536 n460 n378 VDD VSS MUX2_X1 
XU379 n1604 n376 n487 n377 VDD VSS MUX2_X1 
XU378 n1597 n1593 n460 n376 VDD VSS MUX2_X1 
XU377 n375 n357 addr[6] d[8] VDD VSS MUX2_X1 
XU723 n1501 n537 n445 n709 VDD VSS MUX2_X1 
XU722 n708 n696 n433 d[11] VDD VSS MUX2_X1 
XU721 n707 n700 n439 n708 VDD VSS MUX2_X1 
XU720 n706 n703 n503 n707 VDD VSS MUX2_X1 
XU719 n705 n704 n452 n706 VDD VSS MUX2_X1 
XU718 n604 n538 n473 n705 VDD VSS MUX2_X1 
XU717 n1846 n1776 n462 n704 VDD VSS MUX2_X1 
XU716 n702 n701 n452 n703 VDD VSS MUX2_X1 
XU715 n1528 n493 n473 n702 VDD VSS MUX2_X1 
XU714 n1796 n1833 n473 n701 VDD VSS MUX2_X1 
XU713 n699 n697 n503 n700 VDD VSS MUX2_X1 
XU712 n698 n631 n452 n699 VDD VSS MUX2_X1 
XU711 n1787 n1318 n462 n698 VDD VSS MUX2_X1 
XU710 n630 n574 n452 n697 VDD VSS MUX2_X1 
XU709 n695 n691 n439 n696 VDD VSS MUX2_X1 
XU708 n693 n694 n503 n695 VDD VSS MUX2_X1 
XU706 n1670 n692 n452 n693 VDD VSS MUX2_X1 
XU704 n690 n1663 n503 n691 VDD VSS MUX2_X1 
XU703 n689 n1665 n452 n690 VDD VSS MUX2_X1 
XU701 n688 n673 n433 d[10] VDD VSS MUX2_X1 
XU700 n687 n680 n442 n688 VDD VSS MUX2_X1 
XU699 n686 n683 n503 n687 VDD VSS MUX2_X1 
XU698 n685 n684 n452 n686 VDD VSS MUX2_X1 
XU697 n517 n1774 n473 n685 VDD VSS MUX2_X1 
XU696 n522 n1848 n473 n684 VDD VSS MUX2_X1 
XU695 n682 n681 n452 n683 VDD VSS MUX2_X1 
XU694 n1811 n1333 n473 n682 VDD VSS MUX2_X1 
XU693 n1533 n1775 n475 n681 VDD VSS MUX2_X1 
XU692 n679 n676 n503 n680 VDD VSS MUX2_X1 
XU691 n678 n677 n452 n679 VDD VSS MUX2_X1 
XU690 n629 n533 n473 n678 VDD VSS MUX2_X1 
XU689 n1534 n1789 n473 n677 VDD VSS MUX2_X1 
XU688 n675 n674 n452 n676 VDD VSS MUX2_X1 
XU686 n1318 n535 n473 n674 VDD VSS MUX2_X1 
XU685 n672 n666 n445 n673 VDD VSS MUX2_X1 
XU684 n671 n668 n503 n672 VDD VSS MUX2_X1 
XU683 n670 n669 n452 n671 VDD VSS MUX2_X1 
XU682 n532 n1535 n473 n670 VDD VSS MUX2_X1 
XU681 n1541 n524 n473 n669 VDD VSS MUX2_X1 
XU680 n534 n667 n452 n668 VDD VSS MUX2_X1 
XU679 n536 n513 n473 n667 VDD VSS MUX2_X1 
XU678 n665 n1663 n497 n666 VDD VSS MUX2_X1 
XU676 n1545 n1318 n448 n664 VDD VSS MUX2_X1 
XU675 n663 n648 n433 d[0] VDD VSS MUX2_X1 
XU674 n662 n655 n452 n663 VDD VSS MUX2_X1 
XU673 n661 n658 n497 n662 VDD VSS MUX2_X1 
XU672 n659 n660 n458 n661 VDD VSS MUX2_X1 
XU670 n518 n1544 n443 n659 VDD VSS MUX2_X1 
XU669 n657 n656 n473 n658 VDD VSS MUX2_X1 
XU668 n1822 n1790 n443 n657 VDD VSS MUX2_X1 
XU667 n1526 n1501 n442 n656 VDD VSS MUX2_X1 
XU666 n654 n651 n497 n655 VDD VSS MUX2_X1 
XU665 n653 n652 n473 n654 VDD VSS MUX2_X1 
XU664 n628 n524 n442 n653 VDD VSS MUX2_X1 
XU663 n527 n529 n445 n652 VDD VSS MUX2_X1 
XU662 n650 n649 n473 n651 VDD VSS MUX2_X1 
XU661 n526 n1499 n442 n650 VDD VSS MUX2_X1 
XU660 n1501 n1754 n442 n649 VDD VSS MUX2_X1 
XU659 n647 n640 n452 n648 VDD VSS MUX2_X1 
XU658 n646 n643 n507 n647 VDD VSS MUX2_X1 
XU657 n645 n644 n475 n646 VDD VSS MUX2_X1 
XU656 n1674 n1772 n443 n645 VDD VSS MUX2_X1 
XU655 n1855 n509 n443 n644 VDD VSS MUX2_X1 
XU654 n642 n641 n475 n643 VDD VSS MUX2_X1 
XU653 n521 n1835 n443 n642 VDD VSS MUX2_X1 
XU652 n550 n530 n443 n641 VDD VSS MUX2_X1 
XU651 n639 n636 n503 n640 VDD VSS MUX2_X1 
XU650 n637 n638 n473 n639 VDD VSS MUX2_X1 
XU648 n1773 n1789 n439 n637 VDD VSS MUX2_X1 
XU647 n634 n635 n473 n636 VDD VSS MUX2_X1 
XU645 n1808 n1765 n442 n634 VDD VSS MUX2_X1 
XU644 n517 n464 n633 VDD VSS XOR2_X1 
XU643 n461 n513 n632 VDD VSS XOR2_X1 
XU642 n461 n1538 n631 VDD VSS XOR2_X1 
XU641 n539 n473 n630 VDD VSS XOR2_X1 
XU640 n493 n509 n629 VDD VSS XOR2_X1 
XU639 n520 n513 n628 VDD VSS XOR2_X1 
XU638 n526 n513 n627 VDD VSS XOR2_X1 
XU637 n528 n515 n626 VDD VSS XOR2_X1 
XU634 n512 n1501 n473 n623 VDD VSS MUX2_X1 
XU633 n1318 n480 n509 n622 VDD VSS MUX2_X1 
XU632 n1525 n488 n509 n621 VDD VSS MUX2_X1 
XU631 n1520 n492 n509 n620 VDD VSS MUX2_X1 
XU630 n480 n1318 n513 n619 VDD VSS MUX2_X1 
XU629 n488 n1525 n515 n618 VDD VSS MUX2_X1 
XU628 n493 n1525 n515 n617 VDD VSS MUX2_X1 
XU626 n493 n1522 n509 n615 VDD VSS MUX2_X1 
XU625 n1318 n493 n509 n614 VDD VSS MUX2_X1 
XU624 n528 n492 n515 n613 VDD VSS MUX2_X1 
XU623 n526 n488 n509 n612 VDD VSS MUX2_X1 
XU622 n520 n528 n509 n611 VDD VSS MUX2_X1 
XU621 n533 n520 n509 n610 VDD VSS MUX2_X1 
XU620 n1525 n1520 n509 n609 VDD VSS MUX2_X1 
XU835 n820 n805 n433 d[18] VDD VSS MUX2_X1 
XU834 n819 n812 n455 n820 VDD VSS MUX2_X1 
XU833 n818 n815 n495 n819 VDD VSS MUX2_X1 
XU832 n1756 n816 n458 n818 VDD VSS MUX2_X1 
XU830 n814 n813 n471 n815 VDD VSS MUX2_X1 
XU829 n1838 n1760 n443 n814 VDD VSS MUX2_X1 
XU828 n589 n1543 n443 n813 VDD VSS MUX2_X1 
XU827 n811 n808 n495 n812 VDD VSS MUX2_X1 
XU826 n810 n809 n471 n811 VDD VSS MUX2_X1 
XU825 n1743 n1842 n443 n810 VDD VSS MUX2_X1 
XU824 n531 n1534 n443 n809 VDD VSS MUX2_X1 
XU823 n806 n807 n471 n808 VDD VSS MUX2_X1 
XU821 n532 n572 n443 n806 VDD VSS MUX2_X1 
XU820 n804 n797 n455 n805 VDD VSS MUX2_X1 
XU819 n803 n800 n495 n804 VDD VSS MUX2_X1 
XU818 n802 n801 n471 n803 VDD VSS MUX2_X1 
XU817 n586 n1804 n443 n802 VDD VSS MUX2_X1 
XU816 n1824 n1774 n443 n801 VDD VSS MUX2_X1 
XU815 n799 n798 n471 n800 VDD VSS MUX2_X1 
XU814 n1797 n1760 n443 n799 VDD VSS MUX2_X1 
XU813 n1795 n1535 n443 n798 VDD VSS MUX2_X1 
XU812 n795 n796 n495 n797 VDD VSS MUX2_X1 
XU810 n793 n794 n471 n795 VDD VSS MUX2_X1 
XU808 n1811 n555 n443 n793 VDD VSS MUX2_X1 
XU807 n1500 n539 n458 n792 VDD VSS MUX2_X1 
XU806 n597 n445 n458 n791 VDD VSS MUX2_X1 
XU805 n790 n774 n433 d[17] VDD VSS MUX2_X1 
XU804 n789 n782 n445 n790 VDD VSS MUX2_X1 
XU803 n788 n785 n455 n789 VDD VSS MUX2_X1 
XU802 n787 n786 n495 n788 VDD VSS MUX2_X1 
XU801 n569 n1838 n471 n787 VDD VSS MUX2_X1 
XU800 n1523 n540 n471 n786 VDD VSS MUX2_X1 
XU799 n784 n783 n495 n785 VDD VSS MUX2_X1 
XU798 n1741 n541 n471 n784 VDD VSS MUX2_X1 
XU797 n1742 n1762 n471 n783 VDD VSS MUX2_X1 
XU796 n781 n778 n455 n782 VDD VSS MUX2_X1 
XU795 n780 n779 n495 n781 VDD VSS MUX2_X1 
XU794 n1743 n627 n458 n780 VDD VSS MUX2_X1 
XU793 n1756 n1839 n458 n779 VDD VSS MUX2_X1 
XU792 n777 n775 n495 n778 VDD VSS MUX2_X1 
XU791 n1539 n776 n458 n777 VDD VSS MUX2_X1 
XU789 n1756 n1805 n458 n775 VDD VSS MUX2_X1 
XU788 n773 n766 n445 n774 VDD VSS MUX2_X1 
XU787 n772 n769 n455 n773 VDD VSS MUX2_X1 
XU786 n771 n770 n495 n772 VDD VSS MUX2_X1 
XU785 n1797 n539 n458 n771 VDD VSS MUX2_X1 
XU784 n1756 n573 n458 n770 VDD VSS MUX2_X1 
XU783 n768 n767 n507 n769 VDD VSS MUX2_X1 
XU782 n1761 n1777 n475 n768 VDD VSS MUX2_X1 
XU781 n1744 n1791 n475 n767 VDD VSS MUX2_X1 
XU780 n763 n764 n455 n766 VDD VSS MUX2_X1 
XU778 n762 n761 n495 n763 VDD VSS MUX2_X1 
XU777 n512 n1352 n458 n762 VDD VSS MUX2_X1 
XU776 n760 n1838 n458 n761 VDD VSS MUX2_X1 
XU774 n757 n758 n433 d[14] VDD VSS MUX2_X1 
XU772 n756 n752 n503 n757 VDD VSS MUX2_X1 
XU771 n755 n753 n442 n756 VDD VSS MUX2_X1 
XU770 n754 n632 n452 n755 VDD VSS MUX2_X1 
XU769 n577 n1849 n473 n754 VDD VSS MUX2_X1 
XU768 n513 n1671 n452 n753 VDD VSS MUX2_X1 
XU767 n751 n1663 n445 n752 VDD VSS MUX2_X1 
XU766 n1670 n750 n452 n751 VDD VSS MUX2_X1 
XU764 n749 n737 n433 d[13] VDD VSS MUX2_X1 
XU763 n748 n741 n445 n749 VDD VSS MUX2_X1 
XU762 n747 n744 n448 n748 VDD VSS MUX2_X1 
XU761 n746 n745 n468 n747 VDD VSS MUX2_X1 
XU760 n1832 n577 n497 n746 VDD VSS MUX2_X1 
XU759 n547 n1812 n497 n745 VDD VSS MUX2_X1 
XU758 n743 n742 n468 n744 VDD VSS MUX2_X1 
XU755 n739 n740 n452 n741 VDD VSS MUX2_X1 
XU753 n738 n513 n497 n739 VDD VSS MUX2_X1 
XU752 n581 n1528 n473 n738 VDD VSS MUX2_X1 
XU751 n736 n735 n439 n737 VDD VSS MUX2_X1 
XU749 n733 n732 n448 n735 VDD VSS MUX2_X1 
XU746 n531 n1318 n497 n731 VDD VSS MUX2_X1 
XU745 n730 n715 n433 d[12] VDD VSS MUX2_X1 
XU744 n729 n722 n497 n730 VDD VSS MUX2_X1 
XU743 n728 n725 n455 n729 VDD VSS MUX2_X1 
XU742 n727 n726 n458 n728 VDD VSS MUX2_X1 
XU741 n1763 n1535 n443 n727 VDD VSS MUX2_X1 
XU740 n1839 n628 n445 n726 VDD VSS MUX2_X1 
XU739 n724 n723 n458 n725 VDD VSS MUX2_X1 
XU738 n488 n513 n445 n724 VDD VSS MUX2_X1 
XU737 n535 n539 n445 n723 VDD VSS MUX2_X1 
XU736 n721 n718 n455 n722 VDD VSS MUX2_X1 
XU735 n720 n719 n458 n721 VDD VSS MUX2_X1 
XU734 n569 n536 n445 n720 VDD VSS MUX2_X1 
XU733 n480 n513 n445 n719 VDD VSS MUX2_X1 
XU732 n717 n716 n458 n718 VDD VSS MUX2_X1 
XU730 n531 n516 n445 n716 VDD VSS MUX2_X1 
XU729 n713 n714 n497 n715 VDD VSS MUX2_X1 
XU727 n711 n712 n452 n713 VDD VSS MUX2_X1 
XU725 n710 n709 n468 n711 VDD VSS MUX2_X1 
XU939 n923 n922 n477 n924 VDD VSS MUX2_X1 
XU938 n554 n1545 n500 n923 VDD VSS MUX2_X1 
XU937 n548 n1818 n500 n922 VDD VSS MUX2_X1 
XU936 n920 n913 n439 n921 VDD VSS MUX2_X1 
XU935 n919 n916 n454 n920 VDD VSS MUX2_X1 
XU934 n918 n917 n477 n919 VDD VSS MUX2_X1 
XU933 n563 n760 n507 n918 VDD VSS MUX2_X1 
XU932 n1796 n1815 n499 n917 VDD VSS MUX2_X1 
XU931 n915 n914 n475 n916 VDD VSS MUX2_X1 
XU930 n1853 n1767 n507 n915 VDD VSS MUX2_X1 
XU929 n1520 n548 n507 n914 VDD VSS MUX2_X1 
XU928 n911 n912 n454 n913 VDD VSS MUX2_X1 
XU926 n910 n909 n477 n911 VDD VSS MUX2_X1 
XU924 n1779 n608 n507 n909 VDD VSS MUX2_X1 
XU923 n1542 n523 n499 n908 VDD VSS MUX2_X1 
XU922 n907 n892 n433 d[20] VDD VSS MUX2_X1 
XU921 n906 n900 n443 n907 VDD VSS MUX2_X1 
XU920 n905 n902 n454 n906 VDD VSS MUX2_X1 
XU919 n904 n903 n475 n905 VDD VSS MUX2_X1 
XU918 n1775 n556 n507 n904 VDD VSS MUX2_X1 
XU917 n1785 n1745 n507 n903 VDD VSS MUX2_X1 
XU916 n901 n555 n477 n902 VDD VSS MUX2_X1 
XU915 n557 n488 n499 n901 VDD VSS MUX2_X1 
XU914 n899 n895 n454 n900 VDD VSS MUX2_X1 
XU913 n898 n896 n475 n899 VDD VSS MUX2_X1 
XU912 n517 n897 n507 n898 VDD VSS MUX2_X1 
XU910 n562 n591 n507 n896 VDD VSS MUX2_X1 
XU909 n894 n893 n475 n895 VDD VSS MUX2_X1 
XU908 n1522 n603 n507 n894 VDD VSS MUX2_X1 
XU907 n1789 n1784 n507 n893 VDD VSS MUX2_X1 
XU906 n891 n885 n445 n892 VDD VSS MUX2_X1 
XU905 n890 n888 n455 n891 VDD VSS MUX2_X1 
XU904 n512 n889 n475 n890 VDD VSS MUX2_X1 
XU903 n1333 n523 n507 n889 VDD VSS MUX2_X1 
XU902 n887 n886 n475 n888 VDD VSS MUX2_X1 
XU901 n563 n542 n507 n887 VDD VSS MUX2_X1 
XU900 n1741 n1831 n507 n886 VDD VSS MUX2_X1 
XU899 n882 n883 n448 n885 VDD VSS MUX2_X1 
XU897 n881 n880 n473 n882 VDD VSS MUX2_X1 
XU896 n526 n520 n497 n881 VDD VSS MUX2_X1 
XU895 n527 n538 n507 n880 VDD VSS MUX2_X1 
XU894 n879 n864 n433 d[1] VDD VSS MUX2_X1 
XU893 n878 n871 n439 n879 VDD VSS MUX2_X1 
XU892 n877 n874 n452 n878 VDD VSS MUX2_X1 
XU891 n876 n875 n499 n877 VDD VSS MUX2_X1 
XU890 n1815 n1674 n475 n876 VDD VSS MUX2_X1 
XU889 n1761 n1767 n475 n875 VDD VSS MUX2_X1 
XU888 n872 n873 n503 n874 VDD VSS MUX2_X1 
XU886 n547 n1759 n473 n872 VDD VSS MUX2_X1 
XU885 n870 n867 n452 n871 VDD VSS MUX2_X1 
XU884 n869 n868 n503 n870 VDD VSS MUX2_X1 
XU882 n525 n1853 n475 n868 VDD VSS MUX2_X1 
XU881 n866 n865 n503 n867 VDD VSS MUX2_X1 
XU880 n1759 n1541 n473 n866 VDD VSS MUX2_X1 
XU879 n1520 n581 n473 n865 VDD VSS MUX2_X1 
XU878 n863 n856 n439 n864 VDD VSS MUX2_X1 
XU877 n862 n859 n452 n863 VDD VSS MUX2_X1 
XU876 n861 n860 n503 n862 VDD VSS MUX2_X1 
XU875 n575 n557 n462 n861 VDD VSS MUX2_X1 
XU874 n1778 n1535 n473 n860 VDD VSS MUX2_X1 
XU873 n858 n857 n503 n859 VDD VSS MUX2_X1 
XU872 n515 n410 n462 n858 VDD VSS MUX2_X1 
XU871 n1779 n760 n475 n857 VDD VSS MUX2_X1 
XU870 n853 n854 n452 n856 VDD VSS MUX2_X1 
XU868 n852 n851 n507 n853 VDD VSS MUX2_X1 
XU867 n1525 n1533 n475 n852 VDD VSS MUX2_X1 
XU866 n1674 n1501 n475 n851 VDD VSS MUX2_X1 
XU865 n850 n834 n433 d[19] VDD VSS MUX2_X1 
XU864 n849 n842 n455 n850 VDD VSS MUX2_X1 
XU863 n848 n845 n495 n849 VDD VSS MUX2_X1 
XU862 n847 n846 n458 n848 VDD VSS MUX2_X1 
XU861 n1533 n1521 n443 n847 VDD VSS MUX2_X1 
XU860 n529 n1776 n443 n846 VDD VSS MUX2_X1 
XU859 n843 n844 n458 n845 VDD VSS MUX2_X1 
XU857 n1801 n1817 n443 n843 VDD VSS MUX2_X1 
XU856 n841 n838 n495 n842 VDD VSS MUX2_X1 
XU855 n840 n839 n458 n841 VDD VSS MUX2_X1 
XU854 n1523 n573 n443 n840 VDD VSS MUX2_X1 
XU853 n492 n1530 n445 n839 VDD VSS MUX2_X1 
XU852 n835 n836 n458 n838 VDD VSS MUX2_X1 
XU850 n1545 n1523 n443 n835 VDD VSS MUX2_X1 
XU849 n833 n826 n455 n834 VDD VSS MUX2_X1 
XU848 n832 n829 n495 n833 VDD VSS MUX2_X1 
XU847 n831 n830 n471 n832 VDD VSS MUX2_X1 
XU846 n1754 n1500 n443 n831 VDD VSS MUX2_X1 
XU845 n1850 n1814 n443 n830 VDD VSS MUX2_X1 
XU844 n828 n827 n471 n829 VDD VSS MUX2_X1 
XU843 n1817 n531 n443 n828 VDD VSS MUX2_X1 
XU842 n1808 n1776 n443 n827 VDD VSS MUX2_X1 
XU841 n824 n825 n495 n826 VDD VSS MUX2_X1 
XU839 n822 n823 n458 n824 VDD VSS MUX2_X1 
XU837 n1772 n1781 n443 n822 VDD VSS MUX2_X1 
XU836 n601 n629 n443 n821 VDD VSS MUX2_X1 
XU1039 n1020 n1017 n503 n1021 VDD VSS MUX2_X1 
XU1038 n1019 n1018 n462 n1020 VDD VSS MUX2_X1 
XU1037 n555 n515 n435 n1019 VDD VSS MUX2_X1 
XU1036 n615 n1768 n435 n1018 VDD VSS MUX2_X1 
XU1035 n1016 n1015 n462 n1017 VDD VSS MUX2_X1 
XU1034 n897 n1544 n435 n1016 VDD VSS MUX2_X1 
XU1033 n564 n1746 n435 n1015 VDD VSS MUX2_X1 
XU1032 n1013 n1010 n503 n1014 VDD VSS MUX2_X1 
XU1031 n1012 n1011 n464 n1013 VDD VSS MUX2_X1 
XU1030 n1752 n1747 n435 n1012 VDD VSS MUX2_X1 
XU1029 n1352 n562 n435 n1011 VDD VSS MUX2_X1 
XU1028 n1009 n1008 n462 n1010 VDD VSS MUX2_X1 
XU1027 n593 n617 n435 n1009 VDD VSS MUX2_X1 
XU1026 n537 n493 n435 n1008 VDD VSS MUX2_X1 
XU1025 n1006 n999 n452 n1007 VDD VSS MUX2_X1 
XU1024 n1005 n1002 n507 n1006 VDD VSS MUX2_X1 
XU1023 n1004 n1003 n475 n1005 VDD VSS MUX2_X1 
XU1022 n1756 n584 n435 n1004 VDD VSS MUX2_X1 
XU1021 n566 n629 n435 n1003 VDD VSS MUX2_X1 
XU1020 n1001 n1000 n475 n1002 VDD VSS MUX2_X1 
XU1019 n1840 n1745 n435 n1001 VDD VSS MUX2_X1 
XU1018 n579 n609 n435 n1000 VDD VSS MUX2_X1 
XU1017 n998 n995 n503 n999 VDD VSS MUX2_X1 
XU1016 n996 n997 n462 n998 VDD VSS MUX2_X1 
XU1014 n1755 n615 n435 n996 VDD VSS MUX2_X1 
XU1013 n994 n993 n473 n995 VDD VSS MUX2_X1 
XU1010 n992 n977 n435 d[23] VDD VSS MUX2_X1 
XU1009 n991 n984 n439 n992 VDD VSS MUX2_X1 
XU1008 n990 n987 n454 n991 VDD VSS MUX2_X1 
XU1007 n989 n988 n499 n990 VDD VSS MUX2_X1 
XU1006 n1529 n572 n477 n989 VDD VSS MUX2_X1 
XU1005 n1777 n612 n477 n988 VDD VSS MUX2_X1 
XU1004 n986 n985 n499 n987 VDD VSS MUX2_X1 
XU1003 n571 n1775 n477 n986 VDD VSS MUX2_X1 
XU1002 n1529 n606 n477 n985 VDD VSS MUX2_X1 
XU1001 n983 n980 n454 n984 VDD VSS MUX2_X1 
XU1000 n982 n981 n499 n983 VDD VSS MUX2_X1 
XU999 n492 n586 n477 n982 VDD VSS MUX2_X1 
XU998 n571 n583 n477 n981 VDD VSS MUX2_X1 
XU997 n979 n978 n499 n980 VDD VSS MUX2_X1 
XU996 n1780 n565 n462 n979 VDD VSS MUX2_X1 
XU995 n1783 n602 n462 n978 VDD VSS MUX2_X1 
XU994 n976 n970 n439 n977 VDD VSS MUX2_X1 
XU993 n975 n973 n452 n976 VDD VSS MUX2_X1 
XU992 n547 n974 n428 n975 VDD VSS MUX2_X1 
XU991 n544 n1754 n507 n974 VDD VSS MUX2_X1 
XU990 n972 n971 n507 n973 VDD VSS MUX2_X1 
XU989 n530 n1797 n475 n972 VDD VSS MUX2_X1 
XU988 n1521 n520 n475 n971 VDD VSS MUX2_X1 
XU987 n968 n969 n452 n970 VDD VSS MUX2_X1 
XU985 n967 n966 n503 n968 VDD VSS MUX2_X1 
XU983 n591 n1754 n473 n966 VDD VSS MUX2_X1 
XU982 n1812 n492 n507 n965 VDD VSS MUX2_X1 
XU981 n964 n949 n435 d[22] VDD VSS MUX2_X1 
XU980 n963 n956 n439 n964 VDD VSS MUX2_X1 
XU979 n962 n959 n452 n963 VDD VSS MUX2_X1 
XU978 n961 n960 n507 n962 VDD VSS MUX2_X1 
XU977 n526 n516 n473 n961 VDD VSS MUX2_X1 
XU976 n522 n1743 n475 n960 VDD VSS MUX2_X1 
XU975 n958 n957 n507 n959 VDD VSS MUX2_X1 
XU974 n1799 n1790 n475 n958 VDD VSS MUX2_X1 
XU973 n1541 n595 n475 n957 VDD VSS MUX2_X1 
XU972 n955 n952 n454 n956 VDD VSS MUX2_X1 
XU971 n954 n953 n499 n955 VDD VSS MUX2_X1 
XU970 n1845 n1759 n477 n954 VDD VSS MUX2_X1 
XU969 n1318 n565 n462 n953 VDD VSS MUX2_X1 
XU968 n951 n950 n499 n952 VDD VSS MUX2_X1 
XU967 n1825 n1762 n477 n951 VDD VSS MUX2_X1 
XU966 n527 n588 n477 n950 VDD VSS MUX2_X1 
XU965 n948 n941 n439 n949 VDD VSS MUX2_X1 
XU964 n947 n944 n454 n948 VDD VSS MUX2_X1 
XU963 n946 n945 n499 n947 VDD VSS MUX2_X1 
XU962 n570 n1500 n462 n946 VDD VSS MUX2_X1 
XU961 n776 n564 n462 n945 VDD VSS MUX2_X1 
XU960 n943 n942 n499 n944 VDD VSS MUX2_X1 
XU959 n608 n573 n477 n943 VDD VSS MUX2_X1 
XU958 n1808 n542 n477 n942 VDD VSS MUX2_X1 
XU957 n939 n940 n454 n941 VDD VSS MUX2_X1 
XU955 n938 n937 n499 n939 VDD VSS MUX2_X1 
XU954 n555 n601 n477 n938 VDD VSS MUX2_X1 
XU953 n583 n1787 n477 n937 VDD VSS MUX2_X1 
XU952 n602 n1526 n499 n936 VDD VSS MUX2_X1 
XU951 n935 n921 n435 d[21] VDD VSS MUX2_X1 
XU950 n934 n928 n443 n935 VDD VSS MUX2_X1 
XU949 n933 n930 n452 n934 VDD VSS MUX2_X1 
XU948 n932 n931 n475 n933 VDD VSS MUX2_X1 
XU946 n562 n550 n507 n931 VDD VSS MUX2_X1 
XU945 n929 n1806 n475 n930 VDD VSS MUX2_X1 
XU944 n1760 n583 n507 n929 VDD VSS MUX2_X1 
XU943 n927 n924 n454 n928 VDD VSS MUX2_X1 
XU942 n926 n925 n477 n927 VDD VSS MUX2_X1 
XU941 n410 n517 n499 n926 VDD VSS MUX2_X1 
XU940 n1532 n593 n500 n925 VDD VSS MUX2_X1 
XU1142 n523 n567 n462 n1124 VDD VSS MUX2_X1 
XU1141 n1122 n1119 n452 n1123 VDD VSS MUX2_X1 
XU1140 n1121 n1120 n503 n1122 VDD VSS MUX2_X1 
XU1139 n551 n1543 n473 n1121 VDD VSS MUX2_X1 
XU1138 n1538 n567 n462 n1120 VDD VSS MUX2_X1 
XU1137 n1118 n1667 n503 n1119 VDD VSS MUX2_X1 
XU1136 n539 n1826 n462 n1118 VDD VSS MUX2_X1 
XU1135 n1114 n1115 n439 n1117 VDD VSS MUX2_X1 
XU1133 n1113 n1111 n452 n1114 VDD VSS MUX2_X1 
XU1132 n1112 n623 n503 n1113 VDD VSS MUX2_X1 
XU1130 n1110 n513 n503 n1111 VDD VSS MUX2_X1 
XU1128 n623 n1521 n452 n1109 VDD VSS MUX2_X1 
XU1127 n501 n624 n452 n1108 VDD VSS MUX2_X1 
XU1126 n1107 n1092 n435 d[27] VDD VSS MUX2_X1 
XU1125 n1106 n1099 n439 n1107 VDD VSS MUX2_X1 
XU1124 n1105 n1102 n453 n1106 VDD VSS MUX2_X1 
XU1123 n1104 n1103 n500 n1105 VDD VSS MUX2_X1 
XU1122 n1749 n1825 n464 n1104 VDD VSS MUX2_X1 
XU1121 n565 n545 n464 n1103 VDD VSS MUX2_X1 
XU1120 n1101 n1100 n500 n1102 VDD VSS MUX2_X1 
XU1119 n548 n620 n464 n1101 VDD VSS MUX2_X1 
XU1118 n1841 n1759 n464 n1100 VDD VSS MUX2_X1 
XU1117 n1098 n1095 n452 n1099 VDD VSS MUX2_X1 
XU1116 n1097 n1096 n503 n1098 VDD VSS MUX2_X1 
XU1115 n598 n557 n462 n1097 VDD VSS MUX2_X1 
XU1114 n410 n1805 n462 n1096 VDD VSS MUX2_X1 
XU1113 n1093 n1094 n503 n1095 VDD VSS MUX2_X1 
XU1111 n410 n1826 n462 n1093 VDD VSS MUX2_X1 
XU1110 n1091 n1085 n439 n1092 VDD VSS MUX2_X1 
XU1109 n1090 n1087 n454 n1091 VDD VSS MUX2_X1 
XU1108 n1089 n1088 n499 n1090 VDD VSS MUX2_X1 
XU1107 n1808 n536 n462 n1089 VDD VSS MUX2_X1 
XU1106 n1542 n581 n462 n1088 VDD VSS MUX2_X1 
XU1105 n1538 n1086 n428 n1087 VDD VSS MUX2_X1 
XU1103 n1082 n1083 n454 n1085 VDD VSS MUX2_X1 
XU1101 n1081 n1080 n499 n1082 VDD VSS MUX2_X1 
XU1100 n515 n612 n462 n1081 VDD VSS MUX2_X1 
XU1099 n593 n581 n462 n1080 VDD VSS MUX2_X1 
XU1098 n1079 n1064 n435 d[26] VDD VSS MUX2_X1 
XU1097 n1078 n1071 n439 n1079 VDD VSS MUX2_X1 
XU1096 n1077 n1074 n454 n1078 VDD VSS MUX2_X1 
XU1095 n1076 n1075 n500 n1077 VDD VSS MUX2_X1 
XU1094 n1771 n523 n464 n1076 VDD VSS MUX2_X1 
XU1093 n599 n1333 n464 n1075 VDD VSS MUX2_X1 
XU1092 n1073 n1072 n499 n1074 VDD VSS MUX2_X1 
XU1091 n596 n560 n477 n1073 VDD VSS MUX2_X1 
XU1090 n1742 n1779 n475 n1072 VDD VSS MUX2_X1 
XU1089 n1069 n1067 n454 n1071 VDD VSS MUX2_X1 
XU1088 n1068 n1070 n499 n1069 VDD VSS MUX2_X1 
XU1087 n602 n629 n462 n1068 VDD VSS MUX2_X1 
XU1086 n1066 n1065 n499 n1067 VDD VSS MUX2_X1 
XU1085 n1846 n523 n462 n1066 VDD VSS MUX2_X1 
XU1084 n1748 n619 n462 n1065 VDD VSS MUX2_X1 
XU1083 n1063 n1056 n439 n1064 VDD VSS MUX2_X1 
XU1082 n1062 n1059 n452 n1063 VDD VSS MUX2_X1 
XU1081 n1061 n1060 n503 n1062 VDD VSS MUX2_X1 
XU1079 n1776 n567 n462 n1060 VDD VSS MUX2_X1 
XU1078 n1058 n1057 n499 n1059 VDD VSS MUX2_X1 
XU1077 n566 n1827 n462 n1058 VDD VSS MUX2_X1 
XU1076 n1538 n1541 n462 n1057 VDD VSS MUX2_X1 
XU1075 n1054 n1055 n454 n1056 VDD VSS MUX2_X1 
XU1073 n1053 n1052 n499 n1054 VDD VSS MUX2_X1 
XU1072 IN1 n601 n462 n1053 VDD VSS MUX2_X1 
XU1071 n612 n1833 n462 n1052 VDD VSS MUX2_X1 
XU1070 n536 n628 n499 n1051 VDD VSS MUX2_X1 
XU1069 n1050 n1035 n435 d[25] VDD VSS MUX2_X1 
XU1068 n1049 n1042 n439 n1050 VDD VSS MUX2_X1 
XU1067 n1048 n1045 n452 n1049 VDD VSS MUX2_X1 
XU1066 n1047 n1046 n503 n1048 VDD VSS MUX2_X1 
XU1065 n535 n567 n462 n1047 VDD VSS MUX2_X1 
XU1064 n592 n897 n473 n1046 VDD VSS MUX2_X1 
XU1063 n1044 n1043 n503 n1045 VDD VSS MUX2_X1 
XU1062 n1826 n566 n462 n1044 VDD VSS MUX2_X1 
XU1061 n1805 n598 n462 n1043 VDD VSS MUX2_X1 
XU1060 n1041 n1038 n453 n1042 VDD VSS MUX2_X1 
XU1059 n1040 n1039 n500 n1041 VDD VSS MUX2_X1 
XU1058 n1818 n1795 n475 n1040 VDD VSS MUX2_X1 
XU1057 n1333 n1824 n475 n1039 VDD VSS MUX2_X1 
XU1056 n1037 n1036 n500 n1038 VDD VSS MUX2_X1 
XU1055 n605 n1841 n464 n1037 VDD VSS MUX2_X1 
XU1054 n613 n576 n475 n1036 VDD VSS MUX2_X1 
XU1053 n1034 n1028 n439 n1035 VDD VSS MUX2_X1 
XU1052 n1033 n1031 n454 n1034 VDD VSS MUX2_X1 
XU1051 n1672 n1032 n507 n1033 VDD VSS MUX2_X1 
XU1050 n1839 n573 n475 n1032 VDD VSS MUX2_X1 
XU1049 n1030 n1029 n499 n1031 VDD VSS MUX2_X1 
XU1048 n561 n1789 n462 n1030 VDD VSS MUX2_X1 
XU1047 n557 n533 n462 n1029 VDD VSS MUX2_X1 
XU1046 n1025 n1026 n454 n1028 VDD VSS MUX2_X1 
XU1044 n1024 n1023 n499 n1025 VDD VSS MUX2_X1 
XU1042 n601 n1826 n477 n1023 VDD VSS MUX2_X1 
XU1041 n1022 n1007 n439 d[24] VDD VSS MUX2_X1 
XU1040 n1021 n1014 n452 n1022 VDD VSS MUX2_X1 
XU1248 n1757 n1225 n466 n1226 VDD VSS MUX2_X1 
XU1247 n1318 n614 n502 n1225 VDD VSS MUX2_X1 
XU1246 n1223 n1222 n466 n1224 VDD VSS MUX2_X1 
XU1245 n610 n1772 n502 n1223 VDD VSS MUX2_X1 
XU1244 n528 n570 n500 n1222 VDD VSS MUX2_X1 
XU1243 n1220 n1217 n453 n1221 VDD VSS MUX2_X1 
XU1242 n1219 n1218 n466 n1220 VDD VSS MUX2_X1 
XU1241 n1783 n1532 n502 n1219 VDD VSS MUX2_X1 
XU1240 n625 n1333 n502 n1218 VDD VSS MUX2_X1 
XU1239 n1216 n1215 n466 n1217 VDD VSS MUX2_X1 
XU1238 n1811 n1534 n507 n1216 VDD VSS MUX2_X1 
XU1237 n1791 n606 n502 n1215 VDD VSS MUX2_X1 
XU1236 n1213 n1206 n442 n1214 VDD VSS MUX2_X1 
XU1235 n1212 n1209 n453 n1213 VDD VSS MUX2_X1 
XU1234 n1211 n1210 n466 n1212 VDD VSS MUX2_X1 
XU1233 n610 n615 n502 n1211 VDD VSS MUX2_X1 
XU1232 n1828 n1500 n502 n1210 VDD VSS MUX2_X1 
XU1231 n1208 n1207 n466 n1209 VDD VSS MUX2_X1 
XU1230 n563 n620 n500 n1208 VDD VSS MUX2_X1 
XU1229 n554 n543 n500 n1207 VDD VSS MUX2_X1 
XU1227 n1205 n1202 n453 n1206 VDD VSS MUX2_X1 
XU1226 n1204 n1203 n466 n1205 VDD VSS MUX2_X1 
XU1224 n620 n1763 n502 n1203 VDD VSS MUX2_X1 
XU1223 n1201 n1352 n502 n1202 VDD VSS MUX2_X1 
XU1222 n1791 n1752 n466 n1201 VDD VSS MUX2_X1 
XU1221 n1199 n1200 n433 d[30] VDD VSS MUX2_X1 
XU1219 n1198 n1193 n452 n1199 VDD VSS MUX2_X1 
XU1218 n1197 n1194 n445 n1198 VDD VSS MUX2_X1 
XU1217 n1196 n1195 n503 n1197 VDD VSS MUX2_X1 
XU1216 n615 n565 n473 n1196 VDD VSS MUX2_X1 
XU1215 n776 n1501 n473 n1195 VDD VSS MUX2_X1 
XU1214 n1671 n623 n503 n1194 VDD VSS MUX2_X1 
XU1213 n1191 n1192 n442 n1193 VDD VSS MUX2_X1 
XU1211 n1189 n1190 n503 n1191 VDD VSS MUX2_X1 
XU1209 n512 n1333 n473 n1189 VDD VSS MUX2_X1 
XU1208 n503 n1187 n445 n1188 VDD VSS MUX2_X1 
XU1206 n513 n1185 n452 n1186 VDD VSS MUX2_X1 
XU1205 n1184 n529 n445 n1185 VDD VSS MUX2_X1 
XU1204 n513 n569 n458 n1184 VDD VSS MUX2_X1 
XU1203 n1183 n1169 n433 d[2] VDD VSS MUX2_X1 
XU1202 n1182 n1176 n443 n1183 VDD VSS MUX2_X1 
XU1201 n1181 n1179 n455 n1182 VDD VSS MUX2_X1 
XU1200 n1180 n1806 n458 n1181 VDD VSS MUX2_X1 
XU1199 n606 n1499 n507 n1180 VDD VSS MUX2_X1 
XU1198 n1178 n1177 n458 n1179 VDD VSS MUX2_X1 
XU1197 n1742 n1749 n502 n1178 VDD VSS MUX2_X1 
XU1196 n493 n480 n495 n1177 VDD VSS MUX2_X1 
XU1195 n1175 n1172 n455 n1176 VDD VSS MUX2_X1 
XU1194 n1174 n1173 n471 n1175 VDD VSS MUX2_X1 
XU1193 n604 n583 n507 n1174 VDD VSS MUX2_X1 
XU1192 n1758 n1544 n502 n1173 VDD VSS MUX2_X1 
XU1191 n1170 n1171 n471 n1172 VDD VSS MUX2_X1 
XU1189 n549 n585 n502 n1170 VDD VSS MUX2_X1 
XU1188 n1168 n1161 n443 n1169 VDD VSS MUX2_X1 
XU1187 n1167 n1164 n455 n1168 VDD VSS MUX2_X1 
XU1186 n1165 n1166 n471 n1167 VDD VSS MUX2_X1 
XU1184 n1741 n582 n495 n1165 VDD VSS MUX2_X1 
XU1183 n1163 n1162 n471 n1164 VDD VSS MUX2_X1 
XU1182 n616 n551 n502 n1163 VDD VSS MUX2_X1 
XU1181 n587 n610 n502 n1162 VDD VSS MUX2_X1 
XU1180 n1158 n1159 n455 n1161 VDD VSS MUX2_X1 
XU1178 n1157 n1156 n471 n1158 VDD VSS MUX2_X1 
XU1177 n552 n1752 n502 n1157 VDD VSS MUX2_X1 
XU1176 n625 n1835 n502 n1156 VDD VSS MUX2_X1 
XU1175 n1155 n1141 n442 d[29] VDD VSS MUX2_X1 
XU1174 n1154 n1147 n452 n1155 VDD VSS MUX2_X1 
XU1173 n1153 n1150 n458 n1154 VDD VSS MUX2_X1 
XU1172 n1152 n1151 n495 n1153 VDD VSS MUX2_X1 
XU1171 n1812 n516 n433 n1152 VDD VSS MUX2_X1 
XU1170 n1530 n513 n433 n1151 VDD VSS MUX2_X1 
XU1169 n1149 n1148 n495 n1150 VDD VSS MUX2_X1 
XU1168 n594 n512 n433 n1149 VDD VSS MUX2_X1 
XU1167 n1819 n551 n435 n1148 VDD VSS MUX2_X1 
XU1166 n1146 n1144 n468 n1147 VDD VSS MUX2_X1 
XU1165 n1145 n546 n503 n1146 VDD VSS MUX2_X1 
XU1164 n1542 n512 n433 n1145 VDD VSS MUX2_X1 
XU1163 n1142 n1143 n503 n1144 VDD VSS MUX2_X1 
XU1161 n1832 n1500 n433 n1142 VDD VSS MUX2_X1 
XU1160 n1140 n1135 n452 n1141 VDD VSS MUX2_X1 
XU1159 n1139 n1138 n468 n1140 VDD VSS MUX2_X1 
XU1157 n1136 n1137 n503 n1138 VDD VSS MUX2_X1 
XU1155 n536 n1333 n433 n1136 VDD VSS MUX2_X1 
XU1154 n1134 n1132 n473 n1135 VDD VSS MUX2_X1 
XU1153 n513 n1133 n503 n1134 VDD VSS MUX2_X1 
XU1151 n1585 n431 n503 n1132 VDD VSS MUX2_X1 
XU1150 n1131 n1117 n435 d[28] VDD VSS MUX2_X1 
XU1149 n1130 n1123 n439 n1131 VDD VSS MUX2_X1 
XU1148 n1129 n1126 n452 n1130 VDD VSS MUX2_X1 
XU1147 n1128 n1127 n503 n1129 VDD VSS MUX2_X1 
XU1146 n516 n1768 n462 n1128 VDD VSS MUX2_X1 
XU1145 n533 n606 n462 n1127 VDD VSS MUX2_X1 
XU1144 n1125 n1124 n503 n1126 VDD VSS MUX2_X1 
XU1143 n590 n1789 n462 n1125 VDD VSS MUX2_X1 
XU1352 n1756 n488 n500 n1328 VDD VSS MUX2_X1 
XU1351 n1326 n1323 n453 n1327 VDD VSS MUX2_X1 
XU1350 n1325 n1324 n464 n1326 VDD VSS MUX2_X1 
XU1348 n626 n605 n500 n1324 VDD VSS MUX2_X1 
XU1347 n1321 n1322 n464 n1323 VDD VSS MUX2_X1 
XU1345 n595 n1748 n500 n1321 VDD VSS MUX2_X1 
XU1344 n1320 n1305 n435 d[38] VDD VSS MUX2_X1 
XU1343 n1319 n1312 n442 n1320 VDD VSS MUX2_X1 
XU1342 n13180 n1315 n453 n1319 VDD VSS MUX2_X1 
XU1341 n1317 n1316 n502 n13180 VDD VSS MUX2_X1 
XU1340 n578 n512 n466 n1317 VDD VSS MUX2_X1 
XU1339 n1842 n1799 n466 n1316 VDD VSS MUX2_X1 
XU1338 n1314 n1313 n502 n1315 VDD VSS MUX2_X1 
XU1337 n629 n612 n466 n1314 VDD VSS MUX2_X1 
XU1336 n1822 n584 n466 n1313 VDD VSS MUX2_X1 
XU1335 n1311 n1308 n453 n1312 VDD VSS MUX2_X1 
XU1334 n1309 n1310 n500 n1311 VDD VSS MUX2_X1 
XU1332 n558 n1522 n464 n1309 VDD VSS MUX2_X1 
XU1331 n1306 n1307 n500 n1308 VDD VSS MUX2_X1 
XU1329 n579 n578 n466 n1306 VDD VSS MUX2_X1 
XU1328 n1304 n1297 n442 n1305 VDD VSS MUX2_X1 
XU1327 n1303 n1301 n453 n1304 VDD VSS MUX2_X1 
XU1326 n1672 n1302 n500 n1303 VDD VSS MUX2_X1 
XU1325 n622 n593 n475 n1302 VDD VSS MUX2_X1 
XU1324 n1299 n1298 n500 n1301 VDD VSS MUX2_X1 
XU1322 n1523 n537 n475 n1298 VDD VSS MUX2_X1 
XU1321 n1296 n1292 n453 n1297 VDD VSS MUX2_X1 
XU1320 n1293 n1294 n500 n1296 VDD VSS MUX2_X1 
XU1318 n1766 n1816 n464 n1293 VDD VSS MUX2_X1 
XU1317 n1291 n1290 n500 n1292 VDD VSS MUX2_X1 
XU1315 n1545 n621 n464 n1290 VDD VSS MUX2_X1 
XU1314 n1289 n1274 n435 d[37] VDD VSS MUX2_X1 
XU1313 n1288 n1281 n442 n1289 VDD VSS MUX2_X1 
XU1312 n1287 n1284 n502 n1288 VDD VSS MUX2_X1 
XU1311 n1286 n1285 n466 n1287 VDD VSS MUX2_X1 
XU1309 n1751 n609 n453 n1285 VDD VSS MUX2_X1 
XU1308 n1283 n1282 n466 n1284 VDD VSS MUX2_X1 
XU1307 n579 n1754 n453 n1283 VDD VSS MUX2_X1 
XU1306 n1852 n1855 n453 n1282 VDD VSS MUX2_X1 
XU1305 n1280 n1277 n502 n1281 VDD VSS MUX2_X1 
XU1304 n1279 n1278 n466 n1280 VDD VSS MUX2_X1 
XU1303 n1842 n1832 n453 n1279 VDD VSS MUX2_X1 
XU1302 n493 n552 n453 n1278 VDD VSS MUX2_X1 
XU1301 n1276 n1275 n466 n1277 VDD VSS MUX2_X1 
XU1299 n612 n1758 n453 n1275 VDD VSS MUX2_X1 
XU1298 n1273 n1266 n442 n1274 VDD VSS MUX2_X1 
XU1297 n1272 n1269 n500 n1273 VDD VSS MUX2_X1 
XU1296 n1271 n1270 n464 n1272 VDD VSS MUX2_X1 
XU1295 n1530 n560 n453 n1271 VDD VSS MUX2_X1 
XU1294 n1523 n1828 n453 n1270 VDD VSS MUX2_X1 
XU1293 n1268 n1267 n466 n1269 VDD VSS MUX2_X1 
XU1292 n1742 n520 n453 n1268 VDD VSS MUX2_X1 
XU1291 n1767 n1805 n453 n1267 VDD VSS MUX2_X1 
XU1290 n1265 n1262 n500 n1266 VDD VSS MUX2_X1 
XU1289 n1264 n1263 n466 n1265 VDD VSS MUX2_X1 
XU1288 n1756 n1772 n453 n1264 VDD VSS MUX2_X1 
XU1287 n554 n1543 n453 n1263 VDD VSS MUX2_X1 
XU1286 n1261 n1260 n466 n1262 VDD VSS MUX2_X1 
XU1285 n1827 n625 n453 n1261 VDD VSS MUX2_X1 
XU1284 n1841 n1752 n453 n1260 VDD VSS MUX2_X1 
XU1283 n1259 n1243 n435 d[36] VDD VSS MUX2_X1 
XU1282 n1258 n1250 n443 n1259 VDD VSS MUX2_X1 
XU1281 n1257 n1253 n453 n1258 VDD VSS MUX2_X1 
XU1280 n1256 n1254 n466 n1257 VDD VSS MUX2_X1 
XU1279 n526 n1255 n509 n1256 VDD VSS MUX2_X1 
XU1278 n528 n480 n495 n1255 VDD VSS MUX2_X1 
XU1277 n1835 n559 n502 n1254 VDD VSS MUX2_X1 
XU1276 n1252 n1251 n466 n1253 VDD VSS MUX2_X1 
XU1275 n1852 n611 n502 n1252 VDD VSS MUX2_X1 
XU1274 n612 n1753 n502 n1251 VDD VSS MUX2_X1 
XU1273 n1249 n1246 n453 n1250 VDD VSS MUX2_X1 
XU1272 n1248 n1247 n466 n1249 VDD VSS MUX2_X1 
XU1271 n1805 n603 n502 n1248 VDD VSS MUX2_X1 
XU1270 n1770 n607 n502 n1247 VDD VSS MUX2_X1 
XU1269 n1245 n1244 n466 n1246 VDD VSS MUX2_X1 
XU1268 n1747 n1774 n502 n1245 VDD VSS MUX2_X1 
XU1267 n541 n577 n502 n1244 VDD VSS MUX2_X1 
XU1266 n1242 n1235 n443 n1243 VDD VSS MUX2_X1 
XU1265 n1241 n1238 n453 n1242 VDD VSS MUX2_X1 
XU1264 n1240 n1239 n466 n1241 VDD VSS MUX2_X1 
XU1263 n532 n589 n502 n1240 VDD VSS MUX2_X1 
XU1262 n609 n536 n502 n1239 VDD VSS MUX2_X1 
XU1261 n1237 n1236 n466 n1238 VDD VSS MUX2_X1 
XU1260 n1752 n1797 n502 n1237 VDD VSS MUX2_X1 
XU1259 n1814 n1775 n502 n1236 VDD VSS MUX2_X1 
XU1258 n1234 n1231 n453 n1235 VDD VSS MUX2_X1 
XU1257 n1233 n1232 n466 n1234 VDD VSS MUX2_X1 
XU1256 n1824 n1544 n502 n1233 VDD VSS MUX2_X1 
XU1255 n1826 n610 n502 n1232 VDD VSS MUX2_X1 
XU1254 n1230 n1229 n466 n1231 VDD VSS MUX2_X1 
XU1251 n1228 n1214 n435 d[35] VDD VSS MUX2_X1 
XU1250 n1227 n1221 n442 n1228 VDD VSS MUX2_X1 
XU1249 n1226 n1224 n453 n1227 VDD VSS MUX2_X1 
XU1451 n595 n515 n477 n1426 VDD VSS MUX2_X1 
XU1450 n1761 n601 n477 n1425 VDD VSS MUX2_X1 
XU1449 n1423 n1416 n439 n1424 VDD VSS MUX2_X1 
XU1448 n1422 n1419 n454 n1423 VDD VSS MUX2_X1 
XU1447 n1421 n1420 n500 n1422 VDD VSS MUX2_X1 
XU1446 n1752 n621 n464 n1421 VDD VSS MUX2_X1 
XU1445 n517 n1850 n464 n1420 VDD VSS MUX2_X1 
XU1444 n1418 n1417 n499 n1419 VDD VSS MUX2_X1 
XU1443 n1832 n1761 n477 n1418 VDD VSS MUX2_X1 
XU1442 n515 n590 n477 n1417 VDD VSS MUX2_X1 
XU1441 n1415 n1412 n454 n1416 VDD VSS MUX2_X1 
XU1440 n1414 n1413 n499 n1415 VDD VSS MUX2_X1 
XU1439 n1529 n564 n477 n1414 VDD VSS MUX2_X1 
XU1438 n516 n1530 n477 n1413 VDD VSS MUX2_X1 
XU1437 n1411 n1410 n499 n1412 VDD VSS MUX2_X1 
XU1435 n536 n621 n464 n1410 VDD VSS MUX2_X1 
XU1434 n1409 n1395 n435 d[40] VDD VSS MUX2_X1 
XU1433 n1408 n1402 n442 n1409 VDD VSS MUX2_X1 
XU1432 n1407 n1404 n454 n1408 VDD VSS MUX2_X1 
XU1431 n1406 n1405 n477 n1407 VDD VSS MUX2_X1 
XU1429 n526 n601 n499 n1405 VDD VSS MUX2_X1 
XU1428 n1850 n1403 n428 n1404 VDD VSS MUX2_X1 
XU1427 n1797 n1801 n471 n1403 VDD VSS MUX2_X1 
XU1426 n1401 n1398 n454 n1402 VDD VSS MUX2_X1 
XU1425 n1400 n1399 n477 n1401 VDD VSS MUX2_X1 
XU1424 n608 n1352 n499 n1400 VDD VSS MUX2_X1 
XU1423 n564 n596 n499 n1399 VDD VSS MUX2_X1 
XU1422 n1397 n1396 n477 n1398 VDD VSS MUX2_X1 
XU1421 n611 n581 n499 n1397 VDD VSS MUX2_X1 
XU1420 n526 n1765 n500 n1396 VDD VSS MUX2_X1 
XU1419 n1394 n1387 n442 n1395 VDD VSS MUX2_X1 
XU1418 n1393 n1390 n453 n1394 VDD VSS MUX2_X1 
XU1417 n1392 n1391 n464 n1393 VDD VSS MUX2_X1 
XU1416 n586 n599 n500 n1392 VDD VSS MUX2_X1 
XU1415 n548 n1774 n500 n1391 VDD VSS MUX2_X1 
XU1414 n1389 n1388 n464 n1390 VDD VSS MUX2_X1 
XU1413 n543 n1756 n500 n1389 VDD VSS MUX2_X1 
XU1412 n1771 n1318 n500 n1388 VDD VSS MUX2_X1 
XU1411 n1386 n1383 n453 n1387 VDD VSS MUX2_X1 
XU1410 n1385 n1384 n464 n1386 VDD VSS MUX2_X1 
XU1409 n528 n520 n500 n1385 VDD VSS MUX2_X1 
XU1408 n578 n616 n500 n1384 VDD VSS MUX2_X1 
XU1407 n1382 n1381 n464 n1383 VDD VSS MUX2_X1 
XU1406 n543 n1541 n500 n1382 VDD VSS MUX2_X1 
XU1405 n618 n1352 n500 n1381 VDD VSS MUX2_X1 
XU1404 n1380 n1363 n433 d[3] VDD VSS MUX2_X1 
XU1403 n1379 n1372 n443 n1380 VDD VSS MUX2_X1 
XU1402 n1378 n1375 n453 n1379 VDD VSS MUX2_X1 
XU1401 n1377 n1376 n471 n1378 VDD VSS MUX2_X1 
XU1400 n523 n620 n502 n1377 VDD VSS MUX2_X1 
XU1399 n562 n1776 n502 n1376 VDD VSS MUX2_X1 
XU1398 n1374 n1373 n471 n1375 VDD VSS MUX2_X1 
XU1397 n1539 n1751 n502 n1374 VDD VSS MUX2_X1 
XU1396 n569 n561 n502 n1373 VDD VSS MUX2_X1 
XU1395 n1371 n1367 n453 n1372 VDD VSS MUX2_X1 
XU1394 n1370 n1368 n475 n1371 VDD VSS MUX2_X1 
XU1393 n593 n1369 n502 n1370 VDD VSS MUX2_X1 
XU1391 n1746 n605 n507 n1368 VDD VSS MUX2_X1 
XU1390 n1365 n1364 n471 n1367 VDD VSS MUX2_X1 
XU1388 n1805 n1808 n502 n1364 VDD VSS MUX2_X1 
XU1387 n1362 n1355 n443 n1363 VDD VSS MUX2_X1 
XU1386 n1361 n1358 n453 n1362 VDD VSS MUX2_X1 
XU1385 n1360 n1359 n466 n1361 VDD VSS MUX2_X1 
XU1384 n1814 n550 n502 n1360 VDD VSS MUX2_X1 
XU1383 n1500 n620 n502 n1359 VDD VSS MUX2_X1 
XU1382 n1357 n1356 n475 n1358 VDD VSS MUX2_X1 
XU1381 n1352 n1674 n507 n1357 VDD VSS MUX2_X1 
XU1380 n547 n1746 n507 n1356 VDD VSS MUX2_X1 
XU1379 n13520 n1353 n453 n1355 VDD VSS MUX2_X1 
XU1377 n1351 n1350 n466 n13520 VDD VSS MUX2_X1 
XU1376 n1754 n1745 n502 n1351 VDD VSS MUX2_X1 
XU1375 n611 n1776 n502 n1350 VDD VSS MUX2_X1 
XU1374 n1349 n1335 n435 d[39] VDD VSS MUX2_X1 
XU1373 n1348 n1342 n442 n1349 VDD VSS MUX2_X1 
XU1372 n1347 n1344 n453 n1348 VDD VSS MUX2_X1 
XU1371 n1346 n1345 n466 n1347 VDD VSS MUX2_X1 
XU1370 n598 n540 n500 n1346 VDD VSS MUX2_X1 
XU1369 n1827 n1745 n502 n1345 VDD VSS MUX2_X1 
XU1368 n1757 n1343 n466 n1344 VDD VSS MUX2_X1 
XU1367 n1845 n1826 n500 n1343 VDD VSS MUX2_X1 
XU1366 n1341 n1338 n453 n1342 VDD VSS MUX2_X1 
XU1365 n1340 n1339 n466 n1341 VDD VSS MUX2_X1 
XU1364 n552 n618 n502 n1340 VDD VSS MUX2_X1 
XU1363 n527 n1535 n507 n1339 VDD VSS MUX2_X1 
XU1362 n1337 n1336 n466 n1338 VDD VSS MUX2_X1 
XU1360 n1544 n1796 n502 n1336 VDD VSS MUX2_X1 
XU1359 n1334 n1327 n442 n1335 VDD VSS MUX2_X1 
XU1358 n13330 n1330 n453 n1334 VDD VSS MUX2_X1 
XU1357 n1332 n1331 n464 n13330 VDD VSS MUX2_X1 
XU1356 n625 n529 n500 n1332 VDD VSS MUX2_X1 
XU1355 n570 n1318 n500 n1331 VDD VSS MUX2_X1 
XU1354 n1329 n1328 n464 n1330 VDD VSS MUX2_X1 
XU1353 n1819 n1841 n500 n1329 VDD VSS MUX2_X1 
XU1557 n1520 n488 n509 n1515 VDD VSS MUX2_X1 
XU1556 n1513 n1514 n452 n1116 VDD VSS MUX2_X1 
XU1554 n512 n593 n473 n1513 VDD VSS MUX2_X1 
XU1553 n1525 n1318 n509 n1512 VDD VSS MUX2_X1 
XU1552 n628 n1528 n499 n1084 VDD VSS MUX2_X1 
XU1551 n492 n1760 n475 n1511 VDD VSS MUX2_X1 
XU1550 n560 n1538 n507 n1027 VDD VSS MUX2_X1 
XU1549 n526 n517 n509 n1510 VDD VSS MUX2_X1 
XU1548 n493 n1526 n509 n1509 VDD VSS MUX2_X1 
XU1547 n604 n1535 n507 n1508 VDD VSS MUX2_X1 
XU1546 n492 n488 n515 n1507 VDD VSS MUX2_X1 
XU1545 n1333 n628 n497 n884 VDD VSS MUX2_X1 
XU1544 n1840 n572 n507 n855 VDD VSS MUX2_X1 
XU1543 n526 n493 n509 n1506 VDD VSS MUX2_X1 
XU1542 n488 n1520 n509 n1505 VDD VSS MUX2_X1 
XU1541 n1522 n1816 n507 n765 VDD VSS MUX2_X1 
XU1540 n516 n1543 n473 n1504 VDD VSS MUX2_X1 
XU1539 n513 n525 n468 n734 VDD VSS MUX2_X1 
XU1538 n627 n1501 n473 n1503 VDD VSS MUX2_X1 
XU1537 n513 n1498 n448 n1502 VDD VSS MUX2_X1 
XU1526 n528 n488 n515 n1497 VDD VSS MUX2_X1 
XU1525 n615 n462 n1070 VDD VSS XOR2_X1 
XU1524 n1496 n1482 n435 d[43] VDD VSS MUX2_X1 
XU1523 n1495 n1488 n439 n1496 VDD VSS MUX2_X1 
XU1522 n1494 n1491 n454 n1495 VDD VSS MUX2_X1 
XU1521 n1493 n1492 n499 n1494 VDD VSS MUX2_X1 
XU1520 n1811 n605 n477 n1493 VDD VSS MUX2_X1 
XU1519 n553 n577 n477 n1492 VDD VSS MUX2_X1 
XU1518 n1490 n1489 n499 n1491 VDD VSS MUX2_X1 
XU1517 n563 n1541 n477 n1490 VDD VSS MUX2_X1 
XU1516 n1761 n1533 n477 n1489 VDD VSS MUX2_X1 
XU1515 n1487 n1485 n454 n1488 VDD VSS MUX2_X1 
XU1514 n1673 n1486 n499 n1487 VDD VSS MUX2_X1 
XU1513 n1520 n488 n477 n1486 VDD VSS MUX2_X1 
XU1512 n1484 n1483 n499 n1485 VDD VSS MUX2_X1 
XU1511 n1787 n492 n477 n1484 VDD VSS MUX2_X1 
XU1510 n1542 n564 n477 n1483 VDD VSS MUX2_X1 
XU1509 n1481 n1474 n439 n1482 VDD VSS MUX2_X1 
XU1508 n1480 n1477 n454 n1481 VDD VSS MUX2_X1 
XU1507 n1479 n1478 n499 n1480 VDD VSS MUX2_X1 
XU1506 n1773 IN1 n462 n1479 VDD VSS MUX2_X1 
XU1505 n1755 n612 n462 n1478 VDD VSS MUX2_X1 
XU1504 n1476 n1475 n499 n1477 VDD VSS MUX2_X1 
XU1503 n535 n1318 n462 n1476 VDD VSS MUX2_X1 
XU1502 n516 n567 n462 n1475 VDD VSS MUX2_X1 
XU1501 n1473 n1470 n454 n1474 VDD VSS MUX2_X1 
XU1500 n1472 n1471 n499 n1473 VDD VSS MUX2_X1 
XU1499 n533 n1523 n477 n1472 VDD VSS MUX2_X1 
XU1498 n579 n1533 n477 n1471 VDD VSS MUX2_X1 
XU1497 n1469 n1673 n499 n1470 VDD VSS MUX2_X1 
XU1496 n493 n488 n477 n1469 VDD VSS MUX2_X1 
XU1495 n1468 n1454 n435 d[42] VDD VSS MUX2_X1 
XU1494 n1467 n1460 n442 n1468 VDD VSS MUX2_X1 
XU1493 n1466 n1463 n453 n1467 VDD VSS MUX2_X1 
XU1492 n1465 n1464 n500 n1466 VDD VSS MUX2_X1 
XU1491 n545 n1847 n464 n1465 VDD VSS MUX2_X1 
XU1490 n523 n1852 n464 n1464 VDD VSS MUX2_X1 
XU1489 n1462 n1461 n500 n1463 VDD VSS MUX2_X1 
XU1488 n1832 n593 n464 n1462 VDD VSS MUX2_X1 
XU1487 n1525 n540 n464 n1461 VDD VSS MUX2_X1 
XU1486 n1459 n1457 n453 n1460 VDD VSS MUX2_X1 
XU1485 n1458 n633 n500 n1459 VDD VSS MUX2_X1 
XU1484 n526 n612 n464 n1458 VDD VSS MUX2_X1 
XU1483 n1456 n1455 n500 n1457 VDD VSS MUX2_X1 
XU1482 n1797 n516 n466 n1456 VDD VSS MUX2_X1 
XU1481 n1773 n612 n464 n1455 VDD VSS MUX2_X1 
XU1480 n1453 n1446 n442 n1454 VDD VSS MUX2_X1 
XU1479 n1452 n1449 n454 n1453 VDD VSS MUX2_X1 
XU1478 n1451 n1450 n500 n1452 VDD VSS MUX2_X1 
XU1477 n530 n618 n464 n1451 VDD VSS MUX2_X1 
XU1476 n1844 n1533 n464 n1450 VDD VSS MUX2_X1 
XU1475 n1448 n1447 n500 n1449 VDD VSS MUX2_X1 
XU1473 n516 n530 n477 n1447 VDD VSS MUX2_X1 
XU1472 n1445 n1442 n454 n1446 VDD VSS MUX2_X1 
XU1471 n1444 n1443 n500 n1445 VDD VSS MUX2_X1 
XU1470 n584 n1833 n464 n1444 VDD VSS MUX2_X1 
XU1469 n493 n554 n464 n1443 VDD VSS MUX2_X1 
XU1468 n1441 n1440 n500 n1442 VDD VSS MUX2_X1 
XU1467 n515 n585 n464 n1441 VDD VSS MUX2_X1 
XU1466 n1538 n1543 n464 n1440 VDD VSS MUX2_X1 
XU1465 n1439 n1424 n435 d[41] VDD VSS MUX2_X1 
XU1464 n1438 n1431 n439 n1439 VDD VSS MUX2_X1 
XU1463 n1437 n1434 n454 n1438 VDD VSS MUX2_X1 
XU1462 n1436 n1435 n499 n1437 VDD VSS MUX2_X1 
XU1461 n1545 n605 n477 n1436 VDD VSS MUX2_X1 
XU1460 n531 n1815 n477 n1435 VDD VSS MUX2_X1 
XU1459 n1433 n1432 n499 n1434 VDD VSS MUX2_X1 
XU1458 n1529 n1766 n477 n1433 VDD VSS MUX2_X1 
XU1457 n760 n611 n477 n1432 VDD VSS MUX2_X1 
XU1456 n1430 n1427 n454 n1431 VDD VSS MUX2_X1 
XU1455 n1428 n1429 n499 n1430 VDD VSS MUX2_X1 
XU1453 n535 n575 n477 n1428 VDD VSS MUX2_X1 
XU1452 n1426 n1425 n499 n1427 VDD VSS MUX2_X1 
XU450 n622 n1827 VDD VSS INV_X1 
XU449 n556 n1835 VDD VSS INV_X1 
XU448 n21 n1617 VDD VSS INV_X1 
XU447 n545 n1766 VDD VSS INV_X1 
XU446 n750 n1669 VDD VSS INV_X1 
XU445 n43 n1634 VDD VSS INV_X1 
XU444 n26 n1622 VDD VSS INV_X1 
XU443 n596 n1824 VDD VSS INV_X1 
XU442 n575 n1763 VDD VSS INV_X1 
XU441 n19 n1614 VDD VSS INV_X1 
XU440 n566 n1795 VDD VSS INV_X1 
XU437 n572 n1796 VDD VSS INV_X1 
XU419 n598 n1850 VDD VSS INV_X1 
XU418 n584 n1741 VDD VSS INV_X1 
XU417 n522 n1770 VDD VSS INV_X1 
XU416 n1531 n4 n248 n247 VDD VSS AND3_X1 
XU415 n625 n1758 VDD VSS INV_X1 
XU414 n1522 n1528 n410 VDD VSS NOR2_X1 
XU413 n606 n1779 VDD VSS INV_X1 
XU412 n204 n1650 VDD VSS INV_X1 
XU411 n541 n1767 VDD VSS INV_X1 
XU410 n553 n1674 VDD VSS INV_X1 
XU409 n31 n1625 VDD VSS INV_X1 
XU408 n603 n1759 VDD VSS INV_X1 
XU403 n605 n1778 VDD VSS INV_X1 
XU381 n4 n1610 VDD VSS INV_X1 
XU359 n626 n1844 VDD VSS INV_X1 
XU355 n547 n1833 VDD VSS INV_X1 
XU352 n564 n1775 VDD VSS INV_X1 
XU348 n620 n1841 VDD VSS INV_X1 
XU344 n530 n1771 VDD VSS INV_X1 
XU329 n550 n1790 VDD VSS INV_X1 
XU318 n10 n1646 VDD VSS INV_X1 
XU313 n585 n1742 VDD VSS INV_X1 
XU309 n560 n1808 VDD VSS INV_X1 
XU300 n557 n1789 VDD VSS INV_X1 
XU268 n527 n1811 VDD VSS INV_X1 
XU262 n578 n1832 VDD VSS INV_X1 
XU261 n559 n1765 VDD VSS INV_X1 
XU252 n587 n1743 VDD VSS INV_X1 
XU248 n619 n1826 VDD VSS INV_X1 
XU223 n588 n1805 VDD VSS INV_X1 
XU213 n571 n1776 VDD VSS INV_X1 
XU208 n552 n1754 VDD VSS INV_X1 
XU206 n589 n1797 VDD VSS INV_X1 
XU205 n532 n1791 VDD VSS INV_X1 
XU203 n590 n1761 VDD VSS INV_X1 
XU196 n609 n1745 VDD VSS INV_X1 
XU192 n497 n529 n742 VDD VSS NAND2_X1 
XU191 n502 n1745 n1230 VDD VSS NAND2_X1 
XU170 n1708 n1856 VDD VSS INV_X1 
XU168 n58 n1643 VDD VSS INV_X1 
XU130 n2 n4 n261 VDD VSS NAND2_X1 
XU106 n6 n10 n15 VDD VSS NAND2_X1 
XU58 addr[5] n451 VDD VSS INV_X1 
XU56 n448 n449 VDD VSS INV_X1 
XU55 n6 n4 n48 VDD VSS NAND2_X1 
XU53 n609 n502 n587 n1337 VDD VSS AOI21_X1 
XU44 n443 n444 VDD VSS INV_X1 
XU39 n7 n2 n27 VDD VSS NAND2_X1 
XU37 n519 n1522 n538 VDD VSS NAND2_X1 
XU30 n519 n520 n518 VDD VSS NAND2_X1 
XU22 n543 n1522 n558 VDD VSS NAND2_X1 
XU20 n497 n1701 n1694 VDD VSS NAND2_X1 
XU18 n520 n543 n542 VDD VSS NAND2_X1 
XU13 n9 n10 n8 VDD VSS NAND2_X1 
XU11 addr[7] n437 VDD VSS INV_X1 
XU9 n27 n1607 VDD VSS INV_X1 
XU8 n538 n1755 VDD VSS INV_X1 
XU7 n48 n1611 VDD VSS INV_X1 
XU6 n558 n1773 VDD VSS INV_X1 
XU5 n518 n1756 VDD VSS INV_X1 
XU4 n1688 n408 VDD VSS INV_X1 
XU3 n1664 n408 n409 VDD VSS NAND2_X1 
Xc1_reg_17_ n2059 clk_cts_0 n2022 SYNOPSYS_UNCONNECTED_220 VDD VSS DFF_X1 
XU1564 n629 n593 n462 n1519 VDD VSS MUX2_X1 
XU1563 n520 n528 n502 n1366 VDD VSS MUX2_X1 
XU1562 n1763 n1804 n502 n1354 VDD VSS MUX2_X1 
XU1561 n488 n517 n509 n1518 VDD VSS MUX2_X1 
XU1560 n1538 n1758 n502 n1517 VDD VSS MUX2_X1 
XU1559 n492 n1318 n509 n1516 VDD VSS MUX2_X1 
XU1558 n1505 n1765 n495 n1160 VDD VSS MUX2_X1 
XU543 addr[5] n1540 n46 VDD VSS NAND2_X1 
XU542 n1684 n1589 VDD VSS INV_X1 
XU541 n473 n1521 n750 VDD VSS NAND2_X1 
XU540 n1531 n448 n13 VDD VSS OR2_X1 
XU539 n4 n5 n3 VDD VSS NAND2_X1 
XU538 n531 n528 n582 VDD VSS NAND2_X1 
XU537 addr[7] n55 n248 VDD VSS NAND2_X1 
XU536 n464 n558 n1295 VDD VSS NAND2_X1 
XU535 n526 n543 n776 VDD VSS NAND2_X1 
XU533 addr[5] n2 n58 VDD VSS NAND2_X1 
XU531 n519 n526 n760 VDD VSS NAND2_X1 
XU530 n1701 n1702 n1690 VDD VSS NAND2_X1 
XU529 n448 n1537 n21 VDD VSS NAND2_X1 
XU528 n528 n519 n552 VDD VSS NAND2_X1 
XU527 n509 n1525 n587 VDD VSS NAND2_X1 
XU526 addr[5] n1531 n7 VDD VSS NAND2_X1 
XU525 n522 n528 n530 VDD VSS NAND2_X1 
XU524 addr[5] n1527 n130 VDD VSS NAND2_X1 
XU523 n513 n480 n524 VDD VSS NAND2_X1 
XU522 n6 n448 n19 VDD VSS NAND2_X1 
XU520 n501 IN0 n1685 VDD VSS NOR2_X1 
XU519 n531 n526 n560 VDD VSS NAND2_X1 
XU518 n517 n525 n545 VDD VSS NAND2_X1 
XU517 n517 n531 n541 VDD VSS NAND2_X1 
XU516 n515 n1526 n537 VDD VSS NAND2_X1 
XU515 n480 n513 n1726 VDD VSS NOR2_X1 
XU514 n480 n481 n1693 VDD VSS NOR2_X1 
XU512 n543 n517 n625 VDD VSS NAND2_X1 
XU511 n480 n1524 n1700 VDD VSS NOR2_X1 
XU510 n1589 n1700 n1701 n1676 VDD VSS OAI21_X1 
XU509 n528 n525 n527 VDD VSS NAND2_X1 
XU508 n448 n5 n10 VDD VSS NAND2_X1 
XU507 n521 n520 n548 VDD VSS NAND2_X1 
XU506 n5 n448 n411 VDD VSS XNOR2_X1 
XU505 n517 n522 n523 VDD VSS NAND2_X1 
XU503 n448 n486 n1680 VDD VSS NAND2_X1 
XU502 n513 n1318 n529 VDD VSS NAND2_X1 
XU501 n509 n1522 n522 VDD VSS NAND2_X1 
XU500 n448 n1 n4 VDD VSS NAND2_X1 
XU499 n509 n528 n543 VDD VSS NAND2_X1 
XU496 IN0 n501 n1708 VDD VSS NAND2_X1 
XU495 n509 n517 n519 VDD VSS NAND2_X1 
XU493 n509 n520 n531 VDD VSS NAND2_X1 
XU492 n513 n497 n6 VDD VSS NAND2_X1 
XU490 n533 n525 n532 VDD VSS NAND2_X1 
XU489 n509 n526 n525 VDD VSS NAND2_X1 
XU488 n480 IN0 n1701 VDD VSS NOR2_X1 
XU487 n460 n461 VDD VSS INV_X1 
XU482 addr[0] n501 n2 VDD VSS NAND2_X1 
XU480 n492 n480 n520 VDD VSS NAND2_X1 
XU479 n1680 n1664 VDD VSS INV_X1 
XU478 n39 n1630 VDD VSS INV_X1 
XU477 n18 n1613 VDD VSS INV_X1 
XU476 n1517 n1757 VDD VSS INV_X1 
XU475 n1300 n519 n1307 VDD VSS AND2_X1 
XU474 n607 n1840 VDD VSS INV_X1 
XU473 n34 n1628 VDD VSS INV_X1 
XU472 n24 n1620 VDD VSS INV_X1 
XU471 n50 n1639 VDD VSS INV_X1 
XU470 n47 n1637 VDD VSS INV_X1 
XU469 n20 n1616 VDD VSS INV_X1 
XU468 n221 n1645 VDD VSS INV_X1 
XU467 n613 n1845 VDD VSS INV_X1 
XU466 n3 n1612 VDD VSS INV_X1 
XU465 n611 n1831 VDD VSS INV_X1 
XU464 n610 n1784 VDD VSS INV_X1 
XU463 n56 n1641 VDD VSS INV_X1 
XU462 n32 n1626 VDD VSS INV_X1 
XU461 n22 n1618 VDD VSS INV_X1 
XU460 n591 n1777 VDD VSS INV_X1 
XU459 n595 n1804 VDD VSS INV_X1 
XU458 n570 n1846 VDD VSS INV_X1 
XU457 n1633 n248 n354 VDD VSS NAND2_X1 
XU456 n542 n1836 VDD VSS INV_X1 
XU455 n1836 n1295 n1294 VDD VSS NAND2_X1 
XU454 n51 n1640 VDD VSS INV_X1 
XU453 n582 n1838 VDD VSS INV_X1 
XU452 n49 n1638 VDD VSS INV_X1 
XU451 n576 n1839 VDD VSS INV_X1 
XU1162 n519 n1753 VDD VSS INV_X1 
XU1158 n513 n501 n736 VDD VSS NAND2_X1 
XU1156 n1188 n1186 n1200 VDD VSS NOR2_X1 
XU1152 n220 n223 addr[3] n222 VDD VSS AOI21_X1 
XU1134 n578 n501 n1086 VDD VSS AND2_X1 
XU1131 n443 n517 n844 VDD VSS NOR2_X1 
XU1129 n442 n1547 n638 VDD VSS NOR2_X1 
XU1112 IN0 n1650 n168 VDD VSS NOR2_X1 
XU1104 n585 n507 n627 n1406 VDD VSS AOI21_X1 
XU1102 n1752 n453 n536 n1286 VDD VSS AOI21_X1 
XU1080 n593 n501 n579 n932 VDD VSS OAI21_X1 
XU1074 n608 n1785 VDD VSS INV_X1 
XU1045 n443 n1790 n794 VDD VSS NOR2_X1 
XU1043 n59 n1642 VDD VSS INV_X1 
XU1015 n57 n1644 VDD VSS INV_X1 
XU1012 n13 n1608 VDD VSS INV_X1 
XU1011 n407 n1603 VDD VSS INV_X1 
XU986 n17 n1609 VDD VSS INV_X1 
XU984 n25 n1621 VDD VSS INV_X1 
XU956 n540 n1847 VDD VSS INV_X1 
XU947 n817 n1781 VDD VSS INV_X1 
XU927 n468 n1539 n692 VDD VSS NOR2_X1 
XU925 n452 n534 n694 VDD VSS NOR2_X1 
XU911 n473 n965 n969 VDD VSS NOR2_X1 
XU898 n462 n936 n940 VDD VSS NOR2_X1 
XU887 n521 n526 n1369 VDD VSS NAND2_X1 
XU883 n341 n347 n433 n346 VDD VSS AOI21_X1 
XU869 n1643 n460 n13 n379 VDD VSS AOI21_X1 
XU858 n11 n1591 VDD VSS INV_X1 
XU851 n535 n1295 n1448 VDD VSS NAND2_X1 
XU840 n1116 n1108 n1109 n1115 VDD VSS OAI21_X1 
XU838 n42 n1633 VDD VSS INV_X1 
XU831 n604 n1853 VDD VSS INV_X1 
XU811 n29 n1594 VDD VSS INV_X1 
XU809 n554 n1772 VDD VSS INV_X1 
XU790 n501 n569 n743 VDD VSS NOR2_X1 
XU779 n555 n1855 VDD VSS INV_X1 
XU775 n586 n1762 VDD VSS INV_X1 
XU765 n445 n448 n1687 n1706 VDD VSS OAI21_X1 
XU757 n1706 n1590 VDD VSS INV_X1 
XU756 n38 n1597 VDD VSS INV_X1 
XU754 n35 n1595 VDD VSS INV_X1 
XU750 n41 n1632 VDD VSS INV_X1 
XU748 n8 n1648 VDD VSS INV_X1 
XU747 n402 n403 n401 VDD VSS NAND2_X1 
XU731 n1661 n487 n23 n298 VDD VSS AOI21_X1 
XU728 n55 n1600 VDD VSS INV_X1 
XU726 n1599 n484 n311 n310 VDD VSS AOI21_X1 
XU724 n581 n1849 VDD VSS INV_X1 
XU705 n524 n1849 n501 n1325 VDD VSS OAI21_X1 
XU702 n1510 n1752 VDD VSS INV_X1 
XU687 n416 n1654 VDD VSS INV_X1 
XU677 n44 n1635 VDD VSS INV_X1 
XU671 n415 n1653 VDD VSS INV_X1 
XU649 n419 n1656 VDD VSS INV_X1 
XU646 n418 n1655 VDD VSS INV_X1 
XU636 n414 n1652 VDD VSS INV_X1 
XU635 n1502 n1663 VDD VSS INV_X1 
XU627 n1519 n1673 VDD VSS INV_X1 
XU618 n422 n1659 VDD VSS INV_X1 
XU615 n1511 n1672 VDD VSS INV_X1 
XU611 n1520 n509 n607 VDD VSS NAND2_X1 
XU608 n473 n1499 n1110 VDD VSS NAND2_X1 
XU604 addr[7] n28 n351 VDD VSS NOR2_X1 
XU603 n433 n522 n993 VDD VSS NOR2_X1 
XU598 n442 n1539 n710 VDD VSS NOR2_X1 
XU593 n480 n1524 n198 VDD VSS NOR2_X1 
XU592 n462 n1051 n1055 VDD VSS NOR2_X1 
XU591 n417 n1598 VDD VSS INV_X1 
XU579 n1 n19 n54 VDD VSS NAND2_X1 
XU570 n616 n1783 VDD VSS INV_X1 
XU565 n579 n1812 VDD VSS INV_X1 
XU562 n1524 addr[5] n43 VDD VSS NAND2_X1 
XU561 n1743 n502 n561 n1166 VDD VSS AOI21_X1 
XU560 n1765 n473 n527 n869 VDD VSS AOI21_X1 
XU559 n1816 n477 n571 n1024 VDD VSS AOI21_X1 
XU558 n5 n19 n105 VDD VSS NAND2_X1 
XU555 n471 n472 VDD VSS INV_X1 
XU553 n54 n1615 VDD VSS INV_X1 
XU552 n17 addr[7] n53 n252 VDD VSS AOI21_X1 
XU551 n501 n448 n204 VDD VSS NAND2_X1 
XU550 n1543 n453 n565 n1276 VDD VSS AOI21_X1 
XU549 n1586 n1690 n468 n1689 VDD VSS NAND3_X1 
XU548 n1689 n1687 n1688 n1678 VDD VSS OAI21_X1 
XU547 n464 n563 n1300 VDD VSS NAND2_X1 
XU546 n561 n1774 VDD VSS INV_X1 
XU545 n58 n5 n57 VDD VSS NAND2_X1 
XU544 n1523 n502 n616 n1204 VDD VSS AOI21_X1 
XU1616 n492 n493 VDD VSS INV_X1 
XU1614 n480 n493 n528 VDD VSS NAND2_X1 
XU1613 n488 n493 n526 VDD VSS NAND2_X1 
XU1612 n492 n488 n517 VDD VSS NAND2_X1 
XU1611 n624 n1666 VDD VSS INV_X1 
XU1610 n452 n1666 n1187 VDD VSS NAND2_X1 
XU1609 n1697 addr[0] n1728 VDD VSS AND2_X1 
XU1608 n52 n1599 VDD VSS INV_X1 
XU1607 n484 n1536 n189 VDD VSS NAND2_X1 
XU1606 n1704 n1586 VDD VSS INV_X1 
XU1605 n1680 n1704 n1697 VDD VSS NOR2_X1 
XU1603 n433 n442 n1688 VDD VSS NAND2_X1 
XU1602 n487 n486 n1682 VDD VSS NAND2_X1 
XU1601 n1684 n442 IN0 n1729 VDD VSS OAI21_X1 
XU1600 n448 n442 n1699 VDD VSS NOR2_X1 
XU1598 n487 n488 VDD VSS INV_X2 
XU1589 n30 n1624 VDD VSS INV_X1 
XU1588 n46 n1636 VDD VSS INV_X1 
XU1587 n1508 n1806 VDD VSS INV_X1 
XU1586 n1512 n1749 VDD VSS INV_X1 
XU1585 n420 n1657 VDD VSS INV_X1 
XU1584 n1516 n1828 VDD VSS INV_X1 
XU1583 n1503 n1670 VDD VSS INV_X1 
XU1582 n28 n1623 VDD VSS INV_X1 
XU1581 n412 n1604 VDD VSS INV_X1 
XU1580 n423 n1660 VDD VSS INV_X1 
XU1579 n421 n1658 VDD VSS INV_X1 
XU1578 n425 n1662 VDD VSS INV_X1 
XU1577 n1300 n837 n1299 VDD VSS AND2_X1 
XU1576 n37 n1629 VDD VSS INV_X1 
XU1575 n1505 n1817 VDD VSS INV_X1 
XU1574 n549 n1822 VDD VSS INV_X1 
XU1573 n521 n1768 VDD VSS INV_X1 
XU1572 n1498 n1668 VDD VSS INV_X1 
XU1571 n484 n430 n1540 n317 VDD VSS OAI21_X1 
XU1570 n1635 n317 n316 VDD VSS NAND2_X1 
XU1569 n130 n1649 VDD VSS INV_X1 
XU1568 n621 n1748 VDD VSS INV_X1 
XU1567 n618 n1747 VDD VSS INV_X1 
XU1566 n632 n1667 VDD VSS INV_X1 
XU1565 n615 n1780 VDD VSS INV_X1 
XU1555 n617 n1746 VDD VSS INV_X1 
XU1536 n40 n1631 VDD VSS INV_X1 
XU1535 n599 n1814 VDD VSS INV_X1 
XU1534 n424 n1661 VDD VSS INV_X1 
XU1533 n837 n1842 VDD VSS INV_X1 
XU1532 n602 n1815 VDD VSS INV_X1 
XU1531 n544 n1852 VDD VSS INV_X1 
XU1530 n614 n1825 VDD VSS INV_X1 
XU1529 n592 n1744 VDD VSS INV_X1 
XU1528 n573 n1787 VDD VSS INV_X1 
XU1527 n311 n1605 VDD VSS INV_X1 
XU1474 n36 n1596 VDD VSS INV_X1 
XU1454 n1685 n445 n1683 VDD VSS OR2_X1 
XU1436 n594 n1760 VDD VSS INV_X1 
XU1430 n33 n1627 VDD VSS INV_X1 
XU1392 n463 n731 n732 VDD VSS NOR2_X1 
XU1389 n734 n501 n733 VDD VSS NAND2_X1 
XU1378 n1366 n525 n1365 VDD VSS NAND2_X1 
XU1361 n525 n501 n589 n1171 VDD VSS OAI21_X1 
XU1349 n477 n588 n1411 VDD VSS NAND2_X1 
XU1346 n585 n501 n1322 VDD VSS AND2_X1 
XU1333 n626 n464 n529 n1310 VDD VSS AOI21_X1 
XU1330 n537 n501 n1229 VDD VSS NOR2_X1 
XU1323 n546 n1585 VDD VSS INV_X1 
XU1319 n462 n1543 n1094 VDD VSS NOR2_X1 
XU1316 n1853 n507 n910 VDD VSS NAND2_X1 
XU1310 n462 n908 n912 VDD VSS NOR2_X1 
XU1300 n445 n1541 n635 VDD VSS NOR2_X1 
XU1253 n562 n1848 VDD VSS INV_X1 
XU1252 n448 n1524 n342 VDD VSS NOR2_X1 
XU1228 n2 n10 n328 VDD VSS NAND2_X1 
XU1225 n15 n1647 VDD VSS INV_X1 
XU1220 n7 n1606 VDD VSS INV_X1 
XU1212 n23 n1619 VDD VSS INV_X1 
XU1210 n406 n1602 VDD VSS INV_X1 
XU1207 n435 n1744 n997 VDD VSS NOR2_X1 
XU1190 n600 n821 n825 VDD VSS NOR2_X1 
XU1185 n16 n1593 VDD VSS INV_X1 
XU1179 n1537 n1643 n358 VDD VSS NOR2_X1 
XU1711 n1524 n1729 n472 n434 n1717 VDD VSS NAND4_X1 
XU1710 n1586 n497 n448 n1713 n1716 VDD VSS OAI211_X1 
XU1709 n1716 n1717 n1718 n1719 N13521 VDD VSS NAND4_X1 
XU1708 n1522 n516 n521 VDD VSS OR2_X1 
XU1707 n513 n493 n1686 VDD VSS NOR2_X1 
XU1706 n488 n1686 n1856 n1681 VDD VSS OAI21_X1 
XU1705 n501 n516 n1702 VDD VSS NAND2_X1 
XU1704 n1520 n516 n837 VDD VSS NAND2_X1 
XU1703 n1693 n461 n1687 VDD VSS NAND2_X1 
XU1702 n5 n493 n45 VDD VSS NAND2_X1 
XU1701 n509 n493 n544 VDD VSS NAND2_X1 
XU1700 n577 n628 n444 n717 VDD VSS OAI21_X1 
XU1699 n461 n1762 n444 n600 VDD VSS AOI21_X1 
XU1698 n501 n488 addr[0] n1734 VDD VSS NAND3_X1 
XU1697 n468 n1694 n1734 n1732 VDD VSS AOI21_X1 
XU1696 n2 n451 n29 VDD VSS NAND2_X1 
XU1695 n1522 n516 n817 VDD VSS NAND2_X1 
XU1694 n444 n1690 n468 n1695 VDD VSS AOI21_X1 
XU1693 n1695 n1587 VDD VSS INV_X1 
XU1692 n1587 n468 n1685 n1691 VDD VSS OAI21_X1 
XU1691 n535 n472 n1528 n534 VDD VSS OAI21_X1 
XU1690 addr[0] n449 n311 VDD VSS NAND2_X1 
XU1689 n512 n517 n897 VDD VSS NAND2_X1 
XU1688 n520 n461 n574 VDD VSS NAND2_X1 
XU1687 n512 n433 n488 n1725 VDD VSS OAI21_X1 
XU1686 n1725 n501 n1726 n497 n1723 VDD VSS AOI22_X1 
XU1685 n1524 n451 n36 VDD VSS NAND2_X1 
XU1684 n488 n512 n551 VDD VSS NAND2_X1 
XU1683 n512 n528 n540 VDD VSS NAND2_X1 
XU1682 addr[1] n449 n38 VDD VSS NAND2_X1 
XU1681 n468 n1693 n472 n1694 n1692 VDD VSS OAI22_X1 
XU1680 n480 n512 n581 VDD VSS NAND2_X1 
XU1679 n512 n1526 n539 VDD VSS NAND2_X1 
XU1678 n1676 n1588 VDD VSS INV_X1 
XU1677 n1694 n486 n1698 VDD VSS AND2_X1 
XU1676 n1588 n1697 n1690 n1698 n1699 n1696 VDD VSS AOI221_X1 
XU1675 n1696 n1590 n434 n486 n1684 N4870 VDD VSS OAI221_X1 
XU1674 n1684 n1680 n1681 n1682 n1683 n1679 VDD VSS OAI221_X1 
XU1673 n448 n1691 n1692 n444 n1675 VDD VSS AOI22_X1 
XU1672 n1678 n449 n433 n1679 n1677 VDD VSS AOI22_X1 
XU1671 n1677 n433 n1675 n461 n1676 N5090 VDD VSS OAI221_X1 
XU1670 n501 n1726 n472 n1736 VDD VSS NOR3_X1 
XU1669 n1732 n1586 n1733 n1731 VDD VSS NOR3_X1 
XU1668 n1736 n1735 n461 n1730 VDD VSS AOI21_X1 
XU1667 n1731 n452 n1730 n1664 n434 N13331 VDD VSS OAI221_X1 
XU1666 n520 n512 n569 VDD VSS NAND2_X1 
XU1665 n1318 n512 n535 VDD VSS NAND2_X1 
XU1664 n445 n1680 n1701 n1715 VDD VSS OAI21_X1 
XU1663 addr[0] n1715 n1684 n1714 VDD VSS AOI21_X1 
XU1662 n1714 n1713 n1699 n472 n1589 n1712 VDD VSS AOI221_X1 
XU1661 n492 n512 n555 VDD VSS NAND2_X1 
XU1660 n513 n488 n593 VDD VSS NAND2_X1 
XU1659 n512 n526 n536 VDD VSS NAND2_X1 
XU1658 n526 n1526 VDD VSS INV_X1 
XU1657 n448 n444 n1684 VDD VSS NAND2_X1 
XU1656 n1724 n1722 n1708 n1723 n461 n1720 VDD VSS OAI221_X1 
XU1655 n434 n442 n1524 n1721 VDD VSS NOR3_X1 
XU1654 n1721 n408 n1680 n1699 n1720 n1719 VDD VSS AOI221_X1 
XU1653 n512 n497 n1 VDD VSS NAND2_X1 
XU1652 n533 n512 n616 VDD VSS NAND2_X1 
XU1651 n517 n1525 VDD VSS INV_X1 
XU1650 n501 n516 n5 VDD VSS NAND2_X1 
XU1649 n5 n1524 VDD VSS INV_X1 
XU1648 n583 n1523 VDD VSS INV_X1 
XU1647 n533 n1522 VDD VSS INV_X1 
XU1646 n529 n1521 VDD VSS INV_X1 
XU1645 n528 n1520 VDD VSS INV_X1 
XU1644 n551 n1501 VDD VSS INV_X1 
XU1643 n569 n1500 VDD VSS INV_X1 
XU1642 n535 n1499 VDD VSS INV_X1 
XU1641 n593 n1352 VDD VSS INV_X1 
XU1640 n524 n1333 VDD VSS INV_X1 
XU1639 n520 n1318 VDD VSS INV_X1 
XU1638 n515 n516 VDD VSS INV_X1 
XU1634 addr[0] n512 VDD VSS INV_X2 
XU1623 n500 n501 VDD VSS INV_X2 
XU1804 n12 n1536 VDD VSS INV_X1 
XU1803 n567 n1535 VDD VSS INV_X1 
XU1802 n565 n1534 VDD VSS INV_X1 
XU1801 n563 n1533 VDD VSS INV_X1 
XU1800 n612 n1532 VDD VSS INV_X1 
XU1799 n9 n1531 VDD VSS INV_X1 
XU1798 n629 n1530 VDD VSS INV_X1 
XU1797 n628 n1529 VDD VSS INV_X1 
XU1796 n531 n1528 VDD VSS INV_X1 
XU1795 n2 n1527 VDD VSS INV_X1 
XU1794 n45 n1851 VDD VSS INV_X1 
XU1793 n12 n493 n166 VDD VSS NAND2_X1 
XU1792 n1515 n1819 VDD VSS INV_X1 
XU1791 n413 n1651 VDD VSS INV_X1 
XU1790 n1506 n1801 VDD VSS INV_X1 
XU1789 n1160 n472 n1159 VDD VSS AND2_X1 
XU1788 n1084 n472 n1083 VDD VSS AND2_X1 
XU1787 n1825 n472 n1291 VDD VSS AND2_X1 
XU1786 n523 n444 n660 VDD VSS AND2_X1 
XU1785 n1501 n434 n1143 VDD VSS NAND2_X1 
XU1784 n513 n434 n431 VDD VSS AND2_X1 
XU1783 n1531 n449 n430 VDD VSS NOR2_X1 
XU1782 n1354 n472 n1353 VDD VSS AND2_X1 
XU1781 n1501 n461 n1190 VDD VSS NAND2_X1 
XU1780 n503 n1669 n1192 VDD VSS NOR2_X1 
XU1779 n1027 n472 n1026 VDD VSS AND2_X1 
XU1778 n884 n461 n883 VDD VSS AND2_X1 
XU1777 n765 n472 n764 VDD VSS AND2_X1 
XU1776 n565 n461 n566 n675 VDD VSS OAI21_X1 
XU1775 n1540 n493 n146 VDD VSS NOR2_X1 
XU1774 n551 n434 n1137 VDD VSS NAND2_X1 
XU1773 n431 n501 n433 n513 n1139 VDD VSS OAI22_X1 
XU1772 n536 n461 n1112 VDD VSS NOR2_X1 
XU1771 n574 n1665 VDD VSS INV_X1 
XU1770 n1545 n461 n689 VDD VSS NOR2_X1 
XU1769 n837 n444 n565 n836 VDD VSS OAI21_X1 
XU1768 n525 n461 n1668 n449 n759 VDD VSS OAI22_X1 
XU1767 n497 n439 n759 n758 VDD VSS AOI21_X1 
XU1766 n513 n445 n714 VDD VSS NOR2_X1 
XU1765 n1538 n497 n580 VDD VSS NOR2_X1 
XU1764 n461 n580 n1500 n501 n740 VDD VSS OAI22_X1 
XU1763 n855 n472 n854 VDD VSS AND2_X1 
XU1762 n551 n1849 n461 n1429 VDD VSS OAI21_X1 
XU1761 n1497 n1816 VDD VSS INV_X1 
XU1760 n488 n492 n429 VDD VSS XNOR2_X1 
XU1759 n548 n444 n597 VDD VSS NOR2_X1 
XU1758 n791 n792 n796 VDD VSS NOR2_X1 
XU1757 n1521 n434 n1133 VDD VSS NOR2_X1 
XU1756 n568 n664 n665 VDD VSS NOR2_X1 
XU1755 n461 n507 n428 VDD VSS XNOR2_X1 
XU1754 n1500 n472 n1498 VDD VSS NAND2_X1 
XU1753 n1687 n449 n448 n1682 n1707 VDD VSS AOI22_X1 
XU1752 n1707 n1688 N4640 VDD VSS NOR2_X1 
XU1751 n201 n444 n200 VDD VSS AND2_X1 
XU1750 n480 n449 n188 VDD VSS NOR2_X1 
XU1749 n434 n547 n546 VDD VSS NAND2_X1 
XU1748 n451 n1527 n16 VDD VSS NAND2_X1 
XU1747 n12 n1646 n488 n193 VDD VSS OAI21_X1 
XU1746 n539 n1778 n434 n994 VDD VSS OAI21_X1 
XU1745 n53 n437 n48 n259 VDD VSS OAI21_X1 
XU1744 n130 n437 n1643 n267 VDD VSS OAI21_X1 
XU1743 n817 n444 n1541 n816 VDD VSS OAI21_X1 
XU1742 n1771 n444 n1521 n807 VDD VSS OAI21_X1 
XU1741 n1774 n1534 n461 n1061 VDD VSS OAI21_X1 
XU1740 n36 n13 n488 n211 VDD VSS OAI21_X1 
XU1739 n593 n1501 n472 n873 VDD VSS OAI21_X1 
XU1738 n1783 n472 n1543 n967 VDD VSS OAI21_X1 
XU1737 n62 n1601 VDD VSS INV_X1 
XU1736 n130 n488 n1601 n129 VDD VSS OAI21_X1 
XU1735 n1499 n472 n1514 VDD VSS NAND2_X1 
XU1734 n1518 n1751 VDD VSS INV_X1 
XU1733 n1509 n1799 VDD VSS INV_X1 
XU1732 n1504 n1671 VDD VSS INV_X1 
XU1731 n1507 n1818 VDD VSS INV_X1 
XU1730 n6 n449 n427 VDD VSS AND2_X1 
XU1729 n493 n516 n604 VDD VSS NAND2_X1 
XU1728 n460 n21 n426 VDD VSS NAND2_X1 
XU1727 n1525 n516 n592 VDD VSS NAND2_X1 
XU1726 n1 n451 n407 VDD VSS NAND2_X1 
XU1725 n1531 n449 n406 VDD VSS NAND2_X1 
XU1724 n493 n1702 n1705 VDD VSS NOR2_X1 
XU1723 n434 n1664 n1705 n487 n1703 VDD VSS OAI211_X1 
XU1722 n1703 n1704 n1590 n434 N4680 VDD VSS OAI211_X1 
XU1721 n480 n461 n486 n1701 n1711 VDD VSS OAI22_X1 
XU1720 n1712 n497 n1709 VDD VSS OR2_X1 
XU1719 n1699 n497 n1711 n512 n1710 VDD VSS NAND4_X1 
XU1718 n433 n1709 n1710 N19750 VDD VSS AOI21_X1 
XU1717 n449 n1540 n11 VDD VSS NAND2_X1 
XU1716 n1537 n449 n55 VDD VSS NAND2_X1 
XU1715 n29 n484 n11 n306 VDD VSS AOI21_X1 
XU1714 n18 n484 n36 n205 VDD VSS AOI21_X1 
XU1713 n488 n204 n203 VDD VSS NAND2_X1 
XU1712 IN0 n487 n1727 n1728 n1718 VDD VSS OAI211_X1 
XU1849 n445 n472 n520 n712 VDD VSS AND3_X1 
XU1823 n434 n1682 n1699 n1524 N19520 VDD VSS AND4_X1 
XU1822 n444 n488 n38 n207 VDD VSS NAND3_X1 
XU1821 n449 n512 n52 VDD VSS NAND2_X1 
XU1820 n512 n1682 n1713 VDD VSS NAND2_X1 
XU1819 n445 n493 n823 VDD VSS NOR2_X1 
XU1818 n484 n449 n14 VDD VSS NAND2_X1 
XU1817 n497 n472 n624 VDD VSS NAND2_X1 
XU1816 n480 n493 n1524 n1737 VDD VSS NAND3_X1 
XU1815 n1737 n480 n1708 n1735 VDD VSS OAI21_X1 
XU1814 n1684 n1524 n472 n1733 VDD VSS AOI21_X1 
XU1813 n513 n488 n434 n1722 VDD VSS AOI21_X1 
XU1812 n497 n461 n480 n1724 VDD VSS NAND3_X1 
XU1811 n445 n434 n1704 VDD VSS NAND2_X1 
XU1810 n1524 n493 n1740 VDD VSS NAND2_X1 
XU1809 n433 n497 IN0 n480 n1740 n1738 VDD VSS AOI221_X1 
XU1808 n1589 n1586 n1739 VDD VSS NOR2_X1 
XU1807 n1739 n463 n1738 n452 n461 N13181 VDD VSS OAI221_X1 
XU1806 n501 n449 n12 VDD VSS NAND2_X1 
XU1805 n1684 n461 n434 n1727 VDD VSS NOR3_X1 
XCLKBUF_X1_G2B1I1 clk n63_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I3 clk n63_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I4 clk n63_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I5 clk n63_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I7 clk n63_G2B1I7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I9 clk n63_G2B1I9 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I6 clk n63_G2B1I6 VDD VSS CLKBUF_X1 
XU14 n468 n463 VDD VSS BUF_X1 
XU47 d[29] n457 VDD VSS BUF_X1 
XU483 N19750 n459 VDD VSS BUF_X16 
XU485 d[9] n465 VDD VSS INV_X1 
XU494 n465 n467 VDD VSS INV_X32 
XU498 d[8] n469 VDD VSS INV_X1 
XU513 n469 n470 VDD VSS INV_X16 
XU532 d[6] n474 VDD VSS BUF_X1 
XU585 d[5] n476 VDD VSS INV_X1 
XU773 n476 n478 VDD VSS INV_X16 
XU1590 n1856 n479 VDD VSS INV_X1 
XU1592 n479 n481 VDD VSS INV_X8 
XU1593 N4870 n482 VDD VSS INV_X1 
XU1594 n482 n483 VDD VSS INV_X8 
XU1596 n468 n485 VDD VSS INV_X1 
XU1599 n485 n486 VDD VSS INV_X16 
XU1604 N5090 n489 VDD VSS INV_X1 
XU1618 n489 n490 VDD VSS INV_X32 
XU1620 d[48] n491 VDD VSS INV_X1 
XU1626 n491 n494 VDD VSS INV_X32 
XU1627 d[47] n496 VDD VSS BUF_X1 
XU1628 d[46] n498 VDD VSS BUF_X1 
XU1630 d[45] n504 VDD VSS BUF_X1 
XU1632 d[44] n505 VDD VSS INV_X1 
XU1633 n505 n506 VDD VSS INV_X16 
XU1636 N13181 n508 VDD VSS INV_X1 
XU1833 n508 n510 VDD VSS INV_X32 
XU1835 N13331 n511 VDD VSS INV_X1 
XU1836 n511 n514 VDD VSS INV_X32 
XU1837 N13521 n1546 VDD VSS INV_X32 
XU1838 n1546 n1548 VDD VSS INV_X1 
XU1839 n2010 n1549 VDD VSS CLKBUF_X1 
XU1840 n1551 n1550 VDD VSS CLKBUF_X1 
XU1841 n1549 n1551 VDD VSS INV_X32 
XU1842 n1550 c2[16] VDD VSS INV_X32 
XU1843 n2009 n1553 VDD VSS CLKBUF_X1 
XU1844 n1555 n1554 VDD VSS CLKBUF_X1 
XU1845 n1553 n1555 VDD VSS INV_X32 
XU1846 n1554 c2[15] VDD VSS INV_X32 
XU1847 n2008 n1557 VDD VSS CLKBUF_X1 
XU1848 n1559 n1558 VDD VSS CLKBUF_X1 
XU1850 n1557 n1559 VDD VSS INV_X32 
XU1851 n1558 c2[14] VDD VSS INV_X32 
XU1852 n2007 n1561 VDD VSS CLKBUF_X1 
XU1853 n1563 n1562 VDD VSS CLKBUF_X1 
XU1854 n1561 n1563 VDD VSS INV_X32 
XU1855 n1562 c2[13] VDD VSS INV_X32 
XU1856 n2006 n1565 VDD VSS CLKBUF_X1 
XU1857 n1567 n1566 VDD VSS CLKBUF_X1 
XU1858 n1565 n1567 VDD VSS INV_X32 
XU1859 n1566 c2[12] VDD VSS INV_X32 
XU1860 n2018 n1569 VDD VSS CLKBUF_X1 
XU1861 n1571 n1570 VDD VSS CLKBUF_X1 
XU1862 n1569 n1571 VDD VSS INV_X32 
XU1863 n1570 c2[11] VDD VSS INV_X32 
XU1864 n2017 n1573 VDD VSS CLKBUF_X1 
XU1865 n1575 n1574 VDD VSS CLKBUF_X1 
XU1866 n1573 n1575 VDD VSS INV_X32 
XU1867 n1574 c2[10] VDD VSS INV_X32 
XU1868 n2016 n1577 VDD VSS CLKBUF_X1 
XU1869 n1579 n1578 VDD VSS CLKBUF_X1 
XU1870 n1577 n1579 VDD VSS INV_X32 
XU1871 n1578 c2[9] VDD VSS INV_X32 
XU1872 n2015 n1581 VDD VSS CLKBUF_X1 
XU1873 n1583 n1582 VDD VSS CLKBUF_X1 
XU1874 n1581 n1583 VDD VSS INV_X32 
XU1875 n1582 c2[8] VDD VSS INV_X32 
XU1876 n2014 n1592 VDD VSS CLKBUF_X1 
XU1877 n1764 n1750 VDD VSS CLKBUF_X1 
XU1878 n1592 n1764 VDD VSS INV_X32 
XU1879 n1750 c2[7] VDD VSS INV_X32 
XU1880 n2013 n1782 VDD VSS CLKBUF_X1 
XU1881 n1788 n1786 VDD VSS CLKBUF_X1 
XU1882 n1782 n1788 VDD VSS INV_X32 
XU1883 n1786 c2[6] VDD VSS INV_X32 
XU1884 n2012 n1793 VDD VSS CLKBUF_X1 
XU1885 n1798 n1794 VDD VSS CLKBUF_X1 
XU1886 n1793 n1798 VDD VSS INV_X32 
XU1887 n1794 c2[5] VDD VSS INV_X32 
XU1888 n2011 n1802 VDD VSS CLKBUF_X1 
XU1889 n1807 n1803 VDD VSS CLKBUF_X1 
XU1890 n1802 n1807 VDD VSS INV_X32 
XU1891 n1803 c2[4] VDD VSS INV_X32 
XU1892 n2026 n1810 VDD VSS CLKBUF_X1 
XU1893 n1820 n1813 VDD VSS CLKBUF_X1 
XU1894 n1810 n1820 VDD VSS INV_X32 
XU1895 n1813 c2[3] VDD VSS INV_X32 
XU1896 n2025 n1823 VDD VSS CLKBUF_X1 
XU1897 n1830 n1829 VDD VSS CLKBUF_X1 
XU1898 n1823 n1830 VDD VSS INV_X32 
XU1899 n1829 c2[2] VDD VSS INV_X32 
XU1900 n2024 n1837 VDD VSS CLKBUF_X1 
XU1901 n1854 n1843 VDD VSS CLKBUF_X1 
XU1902 n1837 n1854 VDD VSS INV_X32 
XU1903 n1843 c2[1] VDD VSS INV_X32 
XU1904 n2023 n1858 VDD VSS CLKBUF_X1 
XU1905 n1860 n1859 VDD VSS CLKBUF_X1 
XU1906 n1858 n1860 VDD VSS INV_X32 
XU1907 n1859 c2[0] VDD VSS INV_X32 
XU1908 n2058 n1862 VDD VSS CLKBUF_X1 
XU1909 n1864 n1863 VDD VSS CLKBUF_X1 
XU1910 n1862 n1864 VDD VSS INV_X32 
XU1911 n1863 c0[7] VDD VSS INV_X32 
XU1912 n2057 n1866 VDD VSS CLKBUF_X1 
XU1913 n1868 n1867 VDD VSS CLKBUF_X1 
XU1914 n1866 n1868 VDD VSS INV_X32 
XU1915 n1867 c0[6] VDD VSS INV_X32 
XU1916 n2056 n1870 VDD VSS CLKBUF_X1 
XU1917 n1872 n1871 VDD VSS CLKBUF_X1 
XU1918 n1870 n1872 VDD VSS INV_X32 
XU1919 n1871 c0[5] VDD VSS INV_X32 
XU1920 n2055 n1874 VDD VSS CLKBUF_X1 
XU1921 n1876 n1875 VDD VSS CLKBUF_X1 
XU1922 n1874 n1876 VDD VSS INV_X32 
XU1923 n1875 c0[4] VDD VSS INV_X32 
XU1924 n2054 n1878 VDD VSS CLKBUF_X1 
XU1925 n1880 n1879 VDD VSS CLKBUF_X1 
XU1926 n1878 n1880 VDD VSS INV_X32 
XU1927 n1879 c0[3] VDD VSS INV_X32 
XU1928 n2053 n1882 VDD VSS CLKBUF_X1 
XU1929 n1884 n1883 VDD VSS CLKBUF_X1 
XU1930 n1882 n1884 VDD VSS INV_X32 
XU1931 n1883 c0[2] VDD VSS INV_X32 
XU1932 n2052 n1886 VDD VSS CLKBUF_X1 
XU1933 n1888 n1887 VDD VSS CLKBUF_X1 
XU1934 n1886 n1888 VDD VSS INV_X32 
XU1935 n1887 c0[1] VDD VSS INV_X32 
XU1936 n2051 n1890 VDD VSS CLKBUF_X1 
XU1937 n1892 n1891 VDD VSS CLKBUF_X1 
XU1938 n1890 n1892 VDD VSS INV_X32 
XU1939 n1891 c0[0] VDD VSS INV_X32 
XU1940 n2022 n1894 VDD VSS CLKBUF_X1 
XU1941 n1896 n1895 VDD VSS CLKBUF_X1 
XU1942 n1894 n1896 VDD VSS INV_X32 
XU1943 n1895 c1[17] VDD VSS INV_X32 
XU1944 n2021 n1898 VDD VSS CLKBUF_X1 
XU1945 n1900 n1899 VDD VSS CLKBUF_X1 
XU1946 n1898 n1900 VDD VSS INV_X32 
XU1947 n1899 c1[16] VDD VSS INV_X32 
XU1948 n2020 n1902 VDD VSS CLKBUF_X1 
XU1949 n1904 n1903 VDD VSS CLKBUF_X1 
XU1950 n1902 n1904 VDD VSS INV_X32 
XU1951 n1903 c1[15] VDD VSS INV_X32 
XU1952 n2019 n1906 VDD VSS CLKBUF_X1 
XU1953 n1908 n1907 VDD VSS CLKBUF_X1 
XU1954 n1906 n1908 VDD VSS INV_X32 
XU1955 n1907 c1[14] VDD VSS INV_X32 
XU1956 n2034 n1910 VDD VSS CLKBUF_X1 
XU1957 n1912 n1911 VDD VSS CLKBUF_X1 
XU1958 n1910 n1912 VDD VSS INV_X32 
XU1959 n1911 c1[13] VDD VSS INV_X32 
XU1960 n2033 n1914 VDD VSS CLKBUF_X1 
XU1961 n1916 n1915 VDD VSS CLKBUF_X1 
XU1962 n1914 n1916 VDD VSS INV_X32 
XU1963 n1915 c1[12] VDD VSS INV_X32 
XU1964 n1921 c1[11] VDD VSS BUF_X1 
XU1965 n1920 n1919 VDD VSS CLKBUF_X1 
XU1966 n2032 n1920 VDD VSS INV_X32 
XU1967 n1919 n1921 VDD VSS INV_X32 
XU1968 n2031 n1922 VDD VSS CLKBUF_X1 
XU1969 n1924 n1923 VDD VSS CLKBUF_X1 
XU1970 n1922 n1924 VDD VSS INV_X32 
XU1971 n1923 c1[10] VDD VSS INV_X32 
XU1972 n2030 n1926 VDD VSS CLKBUF_X1 
XU1973 n1928 n1927 VDD VSS CLKBUF_X1 
XU1974 n1926 n1928 VDD VSS INV_X32 
XU1975 n1927 c1[9] VDD VSS INV_X32 
XU1976 n2029 n1930 VDD VSS CLKBUF_X1 
XU1977 n1932 n1931 VDD VSS CLKBUF_X1 
XU1978 n1930 n1932 VDD VSS INV_X32 
XU1979 n1931 c1[8] VDD VSS INV_X32 
XU1980 n1937 c1[7] VDD VSS BUF_X1 
XU1981 n1936 n1935 VDD VSS CLKBUF_X1 
XU1982 n2028 n1936 VDD VSS INV_X32 
XU1983 n1935 n1937 VDD VSS INV_X32 
XU1984 n2027 n1938 VDD VSS CLKBUF_X1 
XU1985 n1940 n1939 VDD VSS CLKBUF_X1 
XU1986 n1938 n1940 VDD VSS INV_X32 
XU1987 n1939 c1[6] VDD VSS INV_X32 
XU1988 n2042 n1942 VDD VSS CLKBUF_X1 
XU1989 n1944 n1943 VDD VSS CLKBUF_X1 
XU1990 n1942 n1944 VDD VSS INV_X32 
XU1991 n1943 c1[5] VDD VSS INV_X32 
XU1992 n2041 n1946 VDD VSS CLKBUF_X1 
XU1993 n1948 n1947 VDD VSS CLKBUF_X1 
XU1994 n1946 n1948 VDD VSS INV_X32 
XU1995 n1947 c1[4] VDD VSS INV_X32 
XU1996 n2040 n1950 VDD VSS CLKBUF_X1 
XU1997 n1952 n1951 VDD VSS CLKBUF_X1 
XU1998 n1950 n1952 VDD VSS INV_X32 
XU1999 n1951 c1[3] VDD VSS INV_X32 
XU2000 n1957 c1[2] VDD VSS BUF_X1 
XU2001 n1956 n1955 VDD VSS CLKBUF_X1 
XU2002 n2039 n1956 VDD VSS INV_X32 
XU2003 n1955 n1957 VDD VSS INV_X32 
XU2004 n2038 n1958 VDD VSS CLKBUF_X1 
XU2005 n1960 n1959 VDD VSS CLKBUF_X1 
XU2006 n1958 n1960 VDD VSS INV_X32 
XU2007 n1959 c1[1] VDD VSS INV_X32 
XU2008 n2037 n1962 VDD VSS CLKBUF_X1 
XU2009 n1964 n1963 VDD VSS CLKBUF_X1 
XU2010 n1962 n1964 VDD VSS INV_X32 
XU2011 n1963 c1[0] VDD VSS INV_X32 
XU2012 n2036 n1966 VDD VSS CLKBUF_X1 
XU2013 n1968 n1967 VDD VSS CLKBUF_X1 
XU2014 n1966 n1968 VDD VSS INV_X32 
XU2015 n1967 c0[17] VDD VSS INV_X32 
XU2016 n2035 n1970 VDD VSS CLKBUF_X1 
XU2017 n1972 n1971 VDD VSS CLKBUF_X1 
XU2018 n1970 n1972 VDD VSS INV_X32 
XU2019 n1971 c0[16] VDD VSS INV_X32 
XU2020 n2050 n1974 VDD VSS CLKBUF_X1 
XU2021 n1976 n1975 VDD VSS CLKBUF_X1 
XU2022 n1974 n1976 VDD VSS INV_X32 
XU2023 n1975 c0[15] VDD VSS INV_X32 
XU2024 n2049 n1978 VDD VSS CLKBUF_X1 
XU2025 n1980 n1979 VDD VSS CLKBUF_X1 
XU2026 n1978 n1980 VDD VSS INV_X32 
XU2027 n1979 c0[14] VDD VSS INV_X32 
XU2028 n2048 n1982 VDD VSS CLKBUF_X1 
XU2029 n1984 n1983 VDD VSS CLKBUF_X1 
XU2030 n1982 n1984 VDD VSS INV_X32 
XU2031 n1983 c0[13] VDD VSS INV_X32 
XU2032 n1989 c0[12] VDD VSS BUF_X1 
XU2033 n1988 n1987 VDD VSS CLKBUF_X1 
XU2034 n2047 n1988 VDD VSS INV_X32 
XU2035 n1987 n1989 VDD VSS INV_X32 
XU2036 n2046 n1990 VDD VSS CLKBUF_X1 
XU2037 n1992 n1991 VDD VSS CLKBUF_X1 
XU2038 n1990 n1992 VDD VSS INV_X32 
XU2039 n1991 c0[11] VDD VSS INV_X32 
XU2040 n2045 n1994 VDD VSS CLKBUF_X1 
XU2041 n1996 n1995 VDD VSS CLKBUF_X1 
XU2042 n1994 n1996 VDD VSS INV_X32 
XU2043 n1995 c0[10] VDD VSS INV_X32 
XU2044 n2001 c0[9] VDD VSS BUF_X1 
XU2045 n2000 n1999 VDD VSS CLKBUF_X1 
XU2046 n2044 n2000 VDD VSS INV_X32 
XU2047 n1999 n2001 VDD VSS INV_X32 
XU2048 n2043 n2002 VDD VSS CLKBUF_X1 
XU2049 n2004 n2003 VDD VSS CLKBUF_X1 
XU2050 n2002 n2004 VDD VSS INV_X32 
XU2051 n2003 c0[8] VDD VSS INV_X32 
XU2052 n409 n2059 VDD VSS BUF_X1 
XU2053 n483 n2060 VDD VSS BUF_X1 
XU2054 n510 n2061 VDD VSS BUF_X1 
.ENDS

.SUBCKT gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff clk rstn ce valid_out 
+ VDD VSS IN0 IN1 data_out[63] data_out[62] data_out[61] data_out[60] data_out[59] 
+ data_out[58] data_out[57] data_out[56] data_out[55] data_out[54] data_out[53] 
+ data_out[52] data_out[51] data_out[50] data_out[49] data_out[48] data_out[47] 
+ data_out[46] data_out[45] data_out[44] data_out[43] data_out[42] data_out[41] 
+ data_out[40] data_out[39] data_out[38] data_out[37] data_out[36] data_out[35] 
+ data_out[34] data_out[33] data_out[32] data_out[31] data_out[30] data_out[29] 
+ data_out[28] data_out[27] data_out[26] data_out[25] data_out[24] data_out[23] 
+ data_out[22] data_out[21] data_out[20] data_out[19] data_out[18] data_out[17] 
+ data_out[16] data_out[15] data_out[14] data_out[13] data_out[12] data_out[11] 
+ data_out[10] data_out[9] data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] 
+ data_out[3] data_out[2] data_out[1] data_out[0] IN2 IN3 clk_cts_3 
Xz1_reg_3_ n748 n84_G2B1I5 z1_next[27] n121 VDD VSS DFF_X1 
Xz1_reg_42_ n2007 n78_G2B1I8 z1[42] n79 VDD VSS DFF_X1 
Xz1_reg_18_ n1997 n84 z1_next[42] n106 VDD VSS DFF_X1 
Xz1_reg_52_ n747 n78_G2B1I8 z1[52] n67 VDD VSS DFF_X1 
Xz1_reg_28_ n746 n84_G2B1I3 z1_next[52] n96 VDD VSS DFF_X1 
Xz1_reg_4_ n745 n76_G2B1I4 z1_next[28] n120 VDD VSS DFF_X1 
Xz1_reg_43_ n1976 n84_G2B1I4 z1[43] n77 VDD VSS DFF_X1 
Xz1_reg_19_ n744 n84_G2B1I3 z1_next[43] n105 VDD VSS DFF_X1 
Xz1_reg_53_ n742 n84_G2B1I3 z1[53] n66 VDD VSS DFF_X1 
Xz1_reg_29_ n741 n76_G2B1I4 z1_next[53] n95 VDD VSS DFF_X1 
Xz1_reg_5_ n740 n76_G2B1I4 z1_next[29] n119 VDD VSS DFF_X1 
Xz1_reg_63_ n1949 n84_G2B1I3 SYNOPSYS_UNCONNECTED_643 n56 VDD VSS DFF_X1 
Xz1_reg_39_ n739 n84_G2B1I3 z1_next[63] n85 VDD VSS DFF_X1 
Xz1_reg_15_ n738 n84_G2B1I6 z1_next[39] n109 VDD VSS DFF_X1 
Xz1_reg_49_ n1933 n84_G2B1I6 z1[49] n70 VDD VSS DFF_X1 
Xz1_reg_25_ n734 n84_G2B1I4 z1_next[49] n99 VDD VSS DFF_X1 
Xz1_reg_1_ n1926 n84_G2B1I5 z1_next[25] n123 VDD VSS DFF_X1 
Xz3_reg_61_ n733 n82_G2B1I3 z3[61] n3 VDD VSS DFF_X1 
Xz3_reg_54_ n731 n82_G2B1I7 z3_next[61] n10 VDD VSS DFF_X1 
Xz3_reg_47_ n730 n82_G2B1I3 SYNOPSYS_UNCONNECTED_642 n17 VDD VSS DFF_X1 
Xz3_reg_40_ n728 n80_G2B1I6 SYNOPSYS_UNCONNECTED_641 n24 VDD VSS DFF_X1 
Xz3_reg_33_ n556 n80_G2B1I2 z3_next[40] n31 VDD VSS DFF_X1 
Xz3_reg_26_ n1896 n80_G2B1I6 z3_next[33] n38 VDD VSS DFF_X1 
Xz3_reg_19_ n1891 n80_G2B1I6 SYNOPSYS_UNCONNECTED_640 n45 VDD VSS DFF_X1 
Xz3_reg_12_ n724 n80_G2B1I2 z3_next[19] n52 VDD VSS DFF_X1 
Xz3_reg_57_ n1879 n82_G2B1I3 z3[57] n7 VDD VSS DFF_X1 
Xz3_reg_50_ n722 n82_G2B1I5 SYNOPSYS_UNCONNECTED_639 n14 VDD VSS DFF_X1 
Xz3_reg_43_ n721 n80_G2B1I2 SYNOPSYS_UNCONNECTED_638 n21 VDD VSS DFF_X1 
Xz3_reg_36_ n1861 n76_G2B1I1 z3_next[43] n28 VDD VSS DFF_X1 
Xz3_reg_29_ n720 n76_G2B1I4 z3_next[36] n35 VDD VSS DFF_X1 
Xz3_reg_22_ n718 n76_G2B1I3 SYNOPSYS_UNCONNECTED_637 n42 VDD VSS DFF_X1 
Xz3_reg_15_ n1849 n76_G2B1I3 z3_next[22] n49 VDD VSS DFF_X1 
Xz3_reg_60_ n717 n82_G2B1I4 z3[60] n4 VDD VSS DFF_X1 
Xz3_reg_53_ n1835 n84_G2B1I5 SYNOPSYS_UNCONNECTED_636 n11 VDD VSS DFF_X1 
Xz3_reg_46_ n716 n84_G2B1I5 SYNOPSYS_UNCONNECTED_635 n18 VDD VSS DFF_X1 
Xz3_reg_39_ n715 n84_G2B1I5 z3_next[46] n25 VDD VSS DFF_X1 
Xz3_reg_32_ n714 n84_G2B1I5 z3_next[39] n32 VDD VSS DFF_X1 
Xz3_reg_25_ n713 n80_G2B1I5 z3_next[32] n39 VDD VSS DFF_X1 
Xz3_reg_18_ n712 n84_G2B1I5 SYNOPSYS_UNCONNECTED_634 n46 VDD VSS DFF_X1 
Xz3_reg_11_ n1804 n84_G2B1I2 z3_next[18] n53 VDD VSS DFF_X1 
Xz3_reg_63_ n711 n84_G2B1I4 z3[63] n1 VDD VSS DFF_X1 
Xz3_reg_56_ n710 n82_G2B1I4 z3_next[63] n8 VDD VSS DFF_X1 
Xz3_reg_49_ n1787 clk_G1B1I2 SYNOPSYS_UNCONNECTED_633 n15 VDD VSS DFF_X1 
Xz3_reg_42_ n709 n82_G2B1I8 SYNOPSYS_UNCONNECTED_632 n22 VDD VSS DFF_X1 
Xz3_reg_35_ n708 n82_G2B1I7 z3_next[42] n29 VDD VSS DFF_X1 
Xz3_reg_28_ n1772 n82_G2B1I7 z3_next[35] n36 VDD VSS DFF_X1 
Xz3_reg_21_ n707 n82_G2B1I6 SYNOPSYS_UNCONNECTED_631 n43 VDD VSS DFF_X1 
Xz3_reg_14_ n705 n80_G2B1I6 z3_next[21] n50 VDD VSS DFF_X1 
Xz3_reg_59_ n704 n82_G2B1I3 z3[59] n5 VDD VSS DFF_X1 
Xz3_reg_52_ n702 n82_G2B1I3 SYNOPSYS_UNCONNECTED_630 n12 VDD VSS DFF_X1 
Xz3_reg_45_ n1750 n82_G2B1I6 SYNOPSYS_UNCONNECTED_629 n19 VDD VSS DFF_X1 
Xz3_reg_38_ n1745 n82_G2B1I6 z3_next[45] n26 VDD VSS DFF_X1 
Xz3_reg_31_ n1740 n82_G2B1I5 z3_next[38] n33 VDD VSS DFF_X1 
Xz3_reg_24_ n1731 n76_G2B1I1 z3_next[31] n40 VDD VSS DFF_X1 
Xz3_reg_17_ n697 n76_G2B1I1 z3_next[24] n47 VDD VSS DFF_X1 
Xz3_reg_10_ n1724 n76_G2B1I1 z3_next[17] n54 VDD VSS DFF_X1 
Xz3_reg_62_ n1717 n82_G2B1I3 z3[62] n2 VDD VSS DFF_X1 
Xz3_reg_55_ n695 n82_G2B1I7 z3_next[62] n9 VDD VSS DFF_X1 
Xz3_reg_48_ n1704 n82_G2B1I7 SYNOPSYS_UNCONNECTED_628 n16 VDD VSS DFF_X1 
Xz3_reg_41_ n694 n82_G2B1I7 SYNOPSYS_UNCONNECTED_627 n23 VDD VSS DFF_X1 
Xz3_reg_34_ n693 n82_G2B1I7 z3_next[41] n30 VDD VSS DFF_X1 
Xz3_reg_27_ n1688 n82_G2B1I5 z3_next[34] n37 VDD VSS DFF_X1 
Xz3_reg_20_ n692 n82_G2B1I6 SYNOPSYS_UNCONNECTED_626 n44 VDD VSS DFF_X1 
Xz3_reg_13_ n690 n80_G2B1I6 z3_next[20] n51 VDD VSS DFF_X1 
Xz3_reg_58_ n688 n82_G2B1I7 z3[58] n6 VDD VSS DFF_X1 
Xz3_reg_51_ n687 n82_G2B1I5 z3_next[58] n13 VDD VSS DFF_X1 
Xz3_reg_44_ n686 n82_G2B1I6 SYNOPSYS_UNCONNECTED_625 n20 VDD VSS DFF_X1 
Xz3_reg_37_ n685 n82_G2B1I6 z3_next[44] n27 VDD VSS DFF_X1 
Xz3_reg_30_ n684 n82_G2B1I8 z3_next[37] n34 VDD VSS DFF_X1 
Xz3_reg_23_ n683 n76_G2B1I3 SYNOPSYS_UNCONNECTED_624 n41 VDD VSS DFF_X1 
Xz3_reg_16_ n1644 n76 z3_next[23] n48 VDD VSS DFF_X1 
Xz3_reg_9_ n681 n76_G2B1I1 z3_next[16] n55 VDD VSS DFF_X1 
XU22 n188 n261 VDD VSS BUF_X2 
XU21 n188 n260 VDD VSS BUF_X2 
XU20 n188 n259 VDD VSS BUF_X2 
XU16 n255 n256 VDD VSS INV_X1 
XU12 rstn n252 VDD VSS INV_X1 
XU11 IN0 n250 VDD VSS INV_X1 
XU10 IN1 n248 VDD VSS INV_X1 
XU9 IN3 n246 VDD VSS INV_X1 
XU7 IN2 n185 VDD VSS INV_X1 
Xz2_reg_24_ n1631 n82_G2B1I4 z2_next[37] n166 VDD VSS DFF_X1 
Xz2_reg_11_ n1625 n82_G2B1I4 z2_next[24] n179 VDD VSS DFF_X1 
Xz2_reg_56_ n680 n76_G2B1I1 SYNOPSYS_UNCONNECTED_623 n134 VDD VSS DFF_X1 
Xz2_reg_43_ n679 n76_G2B1I1 z2_next[56] n147 VDD VSS DFF_X1 
Xz2_reg_30_ n678 n76_G2B1I1 z2_next[43] n160 VDD VSS DFF_X1 
Xz2_reg_17_ n1604 n76_G2B1I3 z2_next[30] n173 VDD VSS DFF_X1 
Xz2_reg_62_ n677 n125_G2B1I3 z2[62] n126 VDD VSS DFF_X1 
Xz2_reg_49_ n675 n82_G2B1I8 z2_next[62] n141 VDD VSS DFF_X1 
Xz2_reg_36_ n674 n125_G2B1I3 z2_next[49] n154 VDD VSS DFF_X1 
Xz2_reg_23_ n1587 n76_G2B1I3 z2_next[36] n167 VDD VSS DFF_X1 
Xz2_reg_10_ n1577 n76 z2_next[23] n180 VDD VSS DFF_X1 
Xz2_reg_55_ n672 n125_G2B1I3 SYNOPSYS_UNCONNECTED_622 n135 VDD VSS DFF_X1 
Xz2_reg_42_ n1565 n76 z2_next[55] n148 VDD VSS DFF_X1 
Xz2_reg_29_ n1560 n76_G2B1I4 z2_next[42] n161 VDD VSS DFF_X1 
Xz2_reg_16_ n1554 n76_G2B1I3 z2_next[29] n174 VDD VSS DFF_X1 
Xz2_reg_61_ n671 n125_G2B1I3 z2[61] n128 VDD VSS DFF_X1 
Xz2_reg_48_ n669 n82_G2B1I8 z2_next[61] n142 VDD VSS DFF_X1 
Xz2_reg_35_ n668 n82_G2B1I8 z2_next[48] n155 VDD VSS DFF_X1 
Xz2_reg_22_ n1535 clk_G1B1I2 z2_next[35] n168 VDD VSS DFF_X1 
Xz2_reg_9_ n666 n76_G2B1I1 z2_next[22] n181 VDD VSS DFF_X1 
Xz2_reg_54_ n665 n82_G2B1I8 SYNOPSYS_UNCONNECTED_621 n136 VDD VSS DFF_X1 
Xz2_reg_41_ n663 clk_G1B1I2 z2_next[54] n149 VDD VSS DFF_X1 
Xz2_reg_28_ n662 n82_G2B1I5 z2_next[41] n162 VDD VSS DFF_X1 
Xz2_reg_15_ n661 n82_G2B1I5 z2_next[28] n175 VDD VSS DFF_X1 
Xz2_reg_60_ n659 n82_G2B1I5 SYNOPSYS_UNCONNECTED_620 n130 VDD VSS DFF_X1 
Xz2_reg_47_ n658 n80_G2B1I2 z2_next[60] n143 VDD VSS DFF_X1 
Xz2_reg_34_ n657 n80_G2B1I7 z2_next[47] n156 VDD VSS DFF_X1 
Xz2_reg_21_ n656 n80_G2B1I7 z2_next[34] n169 VDD VSS DFF_X1 
Xz2_reg_8_ n1482 n80_G2B1I7 z2_next[21] n182 VDD VSS DFF_X1 
Xz2_reg_53_ n654 n80_G2B1I4 SYNOPSYS_UNCONNECTED_619 n137 VDD VSS DFF_X1 
Xz2_reg_40_ n653 n80_G2B1I5 z2_next[53] n150 VDD VSS DFF_X1 
Xz2_reg_27_ n651 n80_G2B1I5 z2_next[40] n163 VDD VSS DFF_X1 
Xz2_reg_14_ n1461 n80_G2B1I6 z2_next[27] n176 VDD VSS DFF_X1 
Xz2_reg_59_ n650 n80_G2B1I4 SYNOPSYS_UNCONNECTED_618 n131 VDD VSS DFF_X1 
Xz2_reg_46_ n1450 n80_G2B1I6 z2_next[59] n144 VDD VSS DFF_X1 
Xz2_reg_33_ n649 n80_G2B1I1 z2_next[46] n157 VDD VSS DFF_X1 
Xz2_reg_20_ n1439 n80_G2B1I7 z2_next[33] n170 VDD VSS DFF_X1 
Xz2_reg_7_ n648 n80_G2B1I1 z2_next[20] n183 VDD VSS DFF_X1 
Xz2_reg_52_ n647 n80_G2B1I4 SYNOPSYS_UNCONNECTED_617 n138 VDD VSS DFF_X1 
Xz2_reg_39_ n646 n80_G2B1I2 z2_next[52] n151 VDD VSS DFF_X1 
Xz2_reg_26_ n1422 n80 z2_next[39] n164 VDD VSS DFF_X1 
Xz2_reg_13_ n1412 n80 z2_next[26] n177 VDD VSS DFF_X1 
Xz2_reg_58_ n645 n80_G2B1I4 SYNOPSYS_UNCONNECTED_616 n132 VDD VSS DFF_X1 
Xz2_reg_45_ n642 n80_G2B1I1 z2_next[58] n145 VDD VSS DFF_X1 
Xz2_reg_32_ n1401 n80_G2B1I7 z2_next[45] n158 VDD VSS DFF_X1 
Xz2_reg_19_ n641 n80_G2B1I1 z2_next[32] n171 VDD VSS DFF_X1 
Xz2_reg_6_ n1387 n80_G2B1I5 z2_next[19] n184 VDD VSS DFF_X1 
Xz1_reg_59_ n639 n78_G2B1I7 SYNOPSYS_UNCONNECTED_615 n60 VDD VSS DFF_X1 
Xz1_reg_35_ n638 n80_G2B1I1 z1_next[59] n89 VDD VSS DFF_X1 
Xz1_reg_11_ n636 n78_G2B1I6 z1_next[35] n113 VDD VSS DFF_X1 
Xz1_reg_45_ n635 n78_G2B1I6 z1[45] n74 VDD VSS DFF_X1 
Xz1_reg_21_ n634 n78_G2B1I6 z1_next[45] n103 VDD VSS DFF_X1 
Xz1_reg_60_ n633 n78_G2B1I6 SYNOPSYS_UNCONNECTED_614 n59 VDD VSS DFF_X1 
Xz1_reg_36_ n632 n78_G2B1I7 z1_next[60] n88 VDD VSS DFF_X1 
Xz1_reg_12_ n630 n78_G2B1I4 z1_next[36] n112 VDD VSS DFF_X1 
Xz1_reg_55_ n629 n78_G2B1I2 SYNOPSYS_UNCONNECTED_613 n64 VDD VSS DFF_X1 
Xz1_reg_31_ n628 n84_G2B1I6 z1_next[55] n93 VDD VSS DFF_X1 
Xz1_reg_7_ n627 n84_G2B1I6 z1_next[31] n117 VDD VSS DFF_X1 
Xz1_reg_46_ n617 n78_G2B1I4 z1[46] n73 VDD VSS DFF_X1 
Xz1_reg_22_ n616 n78_G2B1I5 z1_next[46] n102 VDD VSS DFF_X1 
Xz1_reg_61_ n615 n78_G2B1I5 SYNOPSYS_UNCONNECTED_612 n58 VDD VSS DFF_X1 
Xz1_reg_37_ n614 n78_G2B1I2 z1_next[61] n87 VDD VSS DFF_X1 
Xz1_reg_13_ n613 n78_G2B1I4 z1_next[37] n111 VDD VSS DFF_X1 
Xz1_reg_56_ n611 n78_G2B1I8 SYNOPSYS_UNCONNECTED_611 n63 VDD VSS DFF_X1 
Xz1_reg_32_ n608 n78_G2B1I8 z1_next[56] n92 VDD VSS DFF_X1 
Xz1_reg_8_ n1295 n78_G2B1I8 z1_next[32] n116 VDD VSS DFF_X1 
Xz1_reg_47_ n607 n78_G2B1I8 z1[47] n72 VDD VSS DFF_X1 
Xz1_reg_23_ n606 n78_G2B1I5 z1_next[47] n101 VDD VSS DFF_X1 
Xz1_reg_62_ n605 n84 SYNOPSYS_UNCONNECTED_610 n57 VDD VSS DFF_X1 
Xz1_reg_38_ n604 n84_G2B1I4 z1_next[62] n86 VDD VSS DFF_X1 
Xz1_reg_14_ n602 n84_G2B1I6 z1_next[38] n110 VDD VSS DFF_X1 
Xz1_reg_57_ n1261 n78_G2B1I8 SYNOPSYS_UNCONNECTED_609 n62 VDD VSS DFF_X1 
Xz1_reg_33_ n601 n78_G2B1I2 z1_next[57] n91 VDD VSS DFF_X1 
Xz1_reg_9_ n1250 n78_G2B1I2 z1_next[33] n115 VDD VSS DFF_X1 
Xz1_reg_48_ n599 n84_G2B1I4 z1[48] n71 VDD VSS DFF_X1 
Xz1_reg_24_ n598 n76_G2B1I4 z1_next[48] n100 VDD VSS DFF_X1 
Xz1_reg_58_ n1234 n84 SYNOPSYS_UNCONNECTED_608 n61 VDD VSS DFF_X1 
Xz1_reg_34_ n596 n78_G2B1I2 SYNOPSYS_UNCONNECTED_607 n90 VDD VSS DFF_X1 
Xz1_reg_10_ n1228 n78_G2B1I7 z1_next[34] n114 VDD VSS DFF_X1 
Xz1_reg_44_ n594 n84_G2B1I6 z1[44] n75 VDD VSS DFF_X1 
Xz1_reg_20_ n593 n84_G2B1I6 z1_next[44] n104 VDD VSS DFF_X1 
Xz1_reg_54_ n591 n84 z1[54] n65 VDD VSS DFF_X1 
Xz1_reg_30_ n590 n84_G2B1I3 z1_next[54] n94 VDD VSS DFF_X1 
Xz1_reg_6_ n589 n84_G2B1I3 z1_next[30] n118 VDD VSS DFF_X1 
Xz1_reg_40_ n588 n80_G2B1I7 z1[40] n83 VDD VSS DFF_X1 
Xz1_reg_16_ n586 n78_G2B1I6 z1_next[40] n108 VDD VSS DFF_X1 
Xz1_reg_50_ n584 n78_G2B1I7 z1[50] n69 VDD VSS DFF_X1 
Xz1_reg_26_ n583 n80_G2B1I5 z1_next[50] n98 VDD VSS DFF_X1 
Xz1_reg_2_ n582 n80_G2B1I5 z1_next[26] n122 VDD VSS DFF_X1 
Xz1_reg_41_ n1169 n78_G2B1I7 z1[41] n81 VDD VSS DFF_X1 
Xz1_reg_17_ n581 n78_G2B1I6 z1_next[41] n107 VDD VSS DFF_X1 
Xz1_reg_51_ n578 n78_G2B1I4 z1[51] n68 VDD VSS DFF_X1 
Xz1_reg_27_ n577 n84_G2B1I6 z1_next[51] n97 VDD VSS DFF_X1 
XU422 n197 n216 n340 VDD VSS XOR2_X1 
XU421 n231 n340 n339 VDD VSS XOR2_X1 
XU420 n74 z1[50] n215 VDD VSS XOR2_X1 
XU419 n196 n215 n338 VDD VSS XOR2_X1 
XU418 n230 n338 n337 VDD VSS XOR2_X1 
XU417 n73 z1[51] n214 VDD VSS XOR2_X1 
XU416 n195 n214 n336 VDD VSS XOR2_X1 
XU415 n229 n336 n335 VDD VSS XOR2_X1 
XU414 n72 z1[52] n213 VDD VSS XOR2_X1 
XU413 n194 n213 n334 VDD VSS XOR2_X1 
XU412 n228 n334 n333 VDD VSS XOR2_X1 
XU411 n71 z1[53] n212 VDD VSS XOR2_X1 
XU410 n193 n212 n332 VDD VSS XOR2_X1 
XU409 n227 n332 n331 VDD VSS XOR2_X1 
XU408 n70 z1[54] n211 VDD VSS XOR2_X1 
XU407 n192 n211 n330 VDD VSS XOR2_X1 
XU406 n226 n330 n329 VDD VSS XOR2_X1 
Xdata_out_reg_0_ n555 n125_G2B1I6 n2025 SYNOPSYS_UNCONNECTED_606 VDD VSS DFF_X1 
Xdata_out_reg_1_ n1142 n78_G2B1I5 data_out[1] SYNOPSYS_UNCONNECTED_605 VDD VSS DFF_X1 
Xdata_out_reg_2_ n1137 n82_G2B1I3 data_out[2] SYNOPSYS_UNCONNECTED_604 VDD VSS DFF_X1 
Xdata_out_reg_3_ n1132 n82_G2B1I2 data_out[3] SYNOPSYS_UNCONNECTED_603 VDD VSS DFF_X1 
Xdata_out_reg_4_ n1127 n82_G2B1I2 data_out[4] SYNOPSYS_UNCONNECTED_602 VDD VSS DFF_X1 
Xdata_out_reg_5_ n1126 n82_G2B1I2 data_out[5] SYNOPSYS_UNCONNECTED_601 VDD VSS DFF_X1 
Xdata_out_reg_6_ n1118 n82_G2B1I2 n2026 SYNOPSYS_UNCONNECTED_600 VDD VSS DFF_X1 
Xdata_out_reg_7_ n1117 n82_G2B1I7 data_out[7] SYNOPSYS_UNCONNECTED_599 VDD VSS DFF_X1 
Xdata_out_reg_8_ n554 n125_G2B1I5 data_out[8] SYNOPSYS_UNCONNECTED_598 VDD VSS DFF_X1 
Xdata_out_reg_9_ n553 n125_G2B1I5 data_out[9] SYNOPSYS_UNCONNECTED_597 VDD VSS DFF_X1 
Xdata_out_reg_10_ n1098 n82_G2B1I8 data_out[10] SYNOPSYS_UNCONNECTED_596 VDD VSS DFF_X1 
Xdata_out_reg_11_ n1093 n82_G2B1I2 data_out[11] SYNOPSYS_UNCONNECTED_595 VDD VSS DFF_X1 
Xdata_out_reg_12_ n1092 n125 data_out[12] SYNOPSYS_UNCONNECTED_594 VDD VSS DFF_X1 
Xdata_out_reg_13_ n1086 n125 data_out[13] SYNOPSYS_UNCONNECTED_593 VDD VSS DFF_X1 
Xdata_out_reg_14_ n1082 n125 n2024 SYNOPSYS_UNCONNECTED_592 VDD VSS DFF_X1 
Xdata_out_reg_15_ n1076 n125 data_out[15] SYNOPSYS_UNCONNECTED_591 VDD VSS DFF_X1 
Xdata_out_reg_16_ n2028 n125_G2B1I5 data_out[16] SYNOPSYS_UNCONNECTED_590 VDD VSS DFF_X1 
Xdata_out_reg_17_ n1066 n125_G2B1I5 data_out[17] SYNOPSYS_UNCONNECTED_589 VDD VSS DFF_X1 
Xdata_out_reg_18_ n1065 n125_G2B1I1 data_out[18] SYNOPSYS_UNCONNECTED_588 VDD VSS DFF_X1 
Xdata_out_reg_19_ n1056 n125_G2B1I1 data_out[19] SYNOPSYS_UNCONNECTED_587 VDD VSS DFF_X1 
Xdata_out_reg_20_ n1051 n125_G2B1I1 data_out[20] SYNOPSYS_UNCONNECTED_586 VDD VSS DFF_X1 
Xdata_out_reg_21_ n2030 n125_G2B1I3 data_out[21] SYNOPSYS_UNCONNECTED_585 VDD VSS DFF_X1 
Xdata_out_reg_22_ n1044 n125_G2B1I6 data_out[22] SYNOPSYS_UNCONNECTED_584 VDD VSS DFF_X1 
Xdata_out_reg_23_ n1035 n125_G2B1I1 data_out[23] SYNOPSYS_UNCONNECTED_583 VDD VSS DFF_X1 
Xdata_out_reg_24_ n1029 n125_G2B1I6 data_out[24] SYNOPSYS_UNCONNECTED_582 VDD VSS DFF_X1 
Xdata_out_reg_25_ n1023 n76 data_out[25] SYNOPSYS_UNCONNECTED_581 VDD VSS DFF_X1 
Xdata_out_reg_26_ n552 n125_G2B1I3 data_out[26] SYNOPSYS_UNCONNECTED_580 VDD VSS DFF_X1 
Xdata_out_reg_27_ n309 n125_G2B1I1 data_out[27] SYNOPSYS_UNCONNECTED_579 VDD VSS DFF_X1 
Xdata_out_reg_28_ n1009 n76 data_out[28] SYNOPSYS_UNCONNECTED_578 VDD VSS DFF_X1 
Xdata_out_reg_29_ n1003 n125_G2B1I6 data_out[29] SYNOPSYS_UNCONNECTED_577 VDD VSS DFF_X1 
Xdata_out_reg_30_ n997 n125_G2B1I6 data_out[30] SYNOPSYS_UNCONNECTED_576 VDD VSS DFF_X1 
Xdata_out_reg_31_ n308 n125_G2B1I6 data_out[31] SYNOPSYS_UNCONNECTED_575 VDD VSS DFF_X1 
Xdata_out_reg_32_ n985 n78_G2B1I4 data_out[32] SYNOPSYS_UNCONNECTED_574 VDD VSS DFF_X1 
Xdata_out_reg_33_ n979 n78_G2B1I4 data_out[33] SYNOPSYS_UNCONNECTED_573 VDD VSS DFF_X1 
Xdata_out_reg_34_ n973 n78 data_out[34] SYNOPSYS_UNCONNECTED_572 VDD VSS DFF_X1 
Xdata_out_reg_35_ n968 n78_G2B1I6 data_out[35] SYNOPSYS_UNCONNECTED_571 VDD VSS DFF_X1 
Xdata_out_reg_36_ n962 n78_G2B1I1 data_out[36] SYNOPSYS_UNCONNECTED_570 VDD VSS DFF_X1 
Xdata_out_reg_37_ n956 n78_G2B1I1 data_out[37] SYNOPSYS_UNCONNECTED_569 VDD VSS DFF_X1 
Xdata_out_reg_38_ n950 n78_G2B1I5 data_out[38] SYNOPSYS_UNCONNECTED_568 VDD VSS DFF_X1 
Xdata_out_reg_39_ n944 n78_G2B1I4 data_out[39] SYNOPSYS_UNCONNECTED_567 VDD VSS DFF_X1 
Xdata_out_reg_40_ n942 n78 data_out[40] SYNOPSYS_UNCONNECTED_566 VDD VSS DFF_X1 
Xdata_out_reg_41_ n936 n78 data_out[41] SYNOPSYS_UNCONNECTED_565 VDD VSS DFF_X1 
Xdata_out_reg_42_ n573 n78_G2B1I5 data_out[42] SYNOPSYS_UNCONNECTED_564 VDD VSS DFF_X1 
Xdata_out_reg_43_ n924 n78_G2B1I5 data_out[43] SYNOPSYS_UNCONNECTED_563 VDD VSS DFF_X1 
Xdata_out_reg_44_ n918 n78_G2B1I1 data_out[44] SYNOPSYS_UNCONNECTED_562 VDD VSS DFF_X1 
Xdata_out_reg_45_ n307 n78_G2B1I1 data_out[45] SYNOPSYS_UNCONNECTED_561 VDD VSS DFF_X1 
Xdata_out_reg_46_ n906 n78_G2B1I5 data_out[46] SYNOPSYS_UNCONNECTED_560 VDD VSS DFF_X1 
Xdata_out_reg_47_ n900 n78_G2B1I1 data_out[47] SYNOPSYS_UNCONNECTED_559 VDD VSS DFF_X1 
Xdata_out_reg_48_ n894 n125_G2B1I1 data_out[48] SYNOPSYS_UNCONNECTED_558 VDD VSS DFF_X1 
Xdata_out_reg_49_ n888 n125_G2B1I4 data_out[49] SYNOPSYS_UNCONNECTED_557 VDD VSS DFF_X1 
Xdata_out_reg_50_ n882 n125_G2B1I3 data_out[50] SYNOPSYS_UNCONNECTED_556 VDD VSS DFF_X1 
Xdata_out_reg_51_ n306 n125_G2B1I3 data_out[51] SYNOPSYS_UNCONNECTED_555 VDD VSS DFF_X1 
Xdata_out_reg_52_ n870 n125_G2B1I6 data_out[52] SYNOPSYS_UNCONNECTED_554 VDD VSS DFF_X1 
Xdata_out_reg_53_ n864 n125_G2B1I6 data_out[53] SYNOPSYS_UNCONNECTED_553 VDD VSS DFF_X1 
Xdata_out_reg_54_ n858 n125_G2B1I6 data_out[54] SYNOPSYS_UNCONNECTED_552 VDD VSS DFF_X1 
Xdata_out_reg_55_ n852 n125_G2B1I1 data_out[55] SYNOPSYS_UNCONNECTED_551 VDD VSS DFF_X1 
Xdata_out_reg_56_ n846 n125_G2B1I4 data_out[56] SYNOPSYS_UNCONNECTED_550 VDD VSS DFF_X1 
Xdata_out_reg_57_ n305 n125_G2B1I4 data_out[57] SYNOPSYS_UNCONNECTED_549 VDD VSS DFF_X1 
Xdata_out_reg_58_ n836 n125_G2B1I5 data_out[58] SYNOPSYS_UNCONNECTED_548 VDD VSS DFF_X1 
Xdata_out_reg_59_ n2029 n125_G2B1I5 data_out[59] SYNOPSYS_UNCONNECTED_547 VDD VSS DFF_X1 
Xdata_out_reg_60_ n824 n125_G2B1I5 data_out[60] SYNOPSYS_UNCONNECTED_546 VDD VSS DFF_X1 
Xdata_out_reg_61_ n818 n125_G2B1I5 data_out[61] SYNOPSYS_UNCONNECTED_545 VDD VSS DFF_X1 
Xdata_out_reg_62_ n2027 n125_G2B1I4 data_out[62] SYNOPSYS_UNCONNECTED_544 VDD VSS DFF_X1 
Xdata_out_reg_63_ n304 n125_G2B1I4 data_out[63] SYNOPSYS_UNCONNECTED_543 VDD VSS DFF_X1 
Xvalid_out_reg n256 n76_G2B1I3 valid_out SYNOPSYS_UNCONNECTED_542 VDD VSS DFF_X1 
Xz2_reg_51_ n571 n80_G2B1I4 SYNOPSYS_UNCONNECTED_541 n139 VDD VSS DFF_X1 
Xz2_reg_38_ n570 n80_G2B1I6 z2_next[51] n152 VDD VSS DFF_X1 
Xz2_reg_25_ n567 n80 z2_next[38] n165 VDD VSS DFF_X1 
Xz2_reg_12_ n565 n80 z2_next[25] n178 VDD VSS DFF_X1 
Xz2_reg_57_ n564 n80_G2B1I6 SYNOPSYS_UNCONNECTED_540 n133 VDD VSS DFF_X1 
Xz2_reg_44_ n563 n84_G2B1I2 z2_next[57] n146 VDD VSS DFF_X1 
Xz2_reg_31_ n561 n84_G2B1I2 z2_next[44] n159 VDD VSS DFF_X1 
Xz2_reg_18_ n765 n76_G2B1I4 z2_next[31] n172 VDD VSS DFF_X1 
Xz2_reg_63_ n560 n76_G2B1I4 z2[63] n124 VDD VSS DFF_X1 
Xz2_reg_50_ n559 n76_G2B1I1 z2_next[63] n140 VDD VSS DFF_X1 
Xz2_reg_37_ n558 n84_G2B1I2 z2_next[50] n153 VDD VSS DFF_X1 
XU76 IN0 n254 n50 n261 n43 n539 VDD VSS OAI221_X1 
XU75 IN0 n255 n53 n260 n46 n542 VDD VSS OAI221_X1 
XU74 IN0 n254 n729 n261 n24 n520 VDD VSS OAI221_X1 
XU73 IN2 n255 n1646 n258 n41 n537 VDD VSS OAI221_X1 
XU72 IN0 n254 n20 n261 n13 n509 VDD VSS OAI221_X1 
XU71 rstn n254 n13 n261 n1676 n502 VDD VSS OAI221_X1 
XU70 rstn n254 n16 n261 n9 n505 VDD VSS OAI221_X1 
XU69 IN0 n254 n9 n261 n1719 n498 VDD VSS OAI221_X1 
XU68 IN2 n255 n698 n258 n1729 n543 VDD VSS OAI221_X1 
XU67 IN0 n254 n703 n261 n12 n508 VDD VSS OAI221_X1 
XU66 IN0 n254 n12 n261 n5 n501 VDD VSS OAI221_X1 
XU65 rstn n254 n29 n258 n22 n518 VDD VSS OAI221_X1 
XU64 IN2 n255 n22 n258 n1797 n511 VDD VSS OAI221_X1 
XU63 IN0 n254 n1797 n258 n806 n504 VDD VSS OAI221_X1 
XU62 IN2 n255 n806 n260 n1 n497 VDD VSS OAI221_X1 
XU61 IN0 n254 n11 n261 n4 n500 VDD VSS OAI221_X1 
XU60 IN2 n255 n719 n258 n42 n538 VDD VSS OAI221_X1 
XU59 IN0 n254 n14 n261 n1881 n503 VDD VSS OAI221_X1 
XU58 IN0 n254 n1886 n261 n726 n541 VDD VSS OAI221_X1 
XU57 rstn n254 n732 n261 n10 n506 VDD VSS OAI221_X1 
XU56 IN0 n254 n10 n261 n3 n499 VDD VSS OAI221_X1 
XU55 IN3 n2531 n735 n260 n1931 n472 VDD VSS OAI221_X1 
XU54 IN3 n2531 n109 n260 n85 n458 VDD VSS OAI221_X1 
XU53 IN2 n255 n119 n260 n95 n468 VDD VSS OAI221_X1 
XU52 IN2 n255 n120 n260 n96 n469 VDD VSS OAI221_X1 
XU51 IN3 n2531 n96 n259 n67 n445 VDD VSS OAI221_X1 
XU50 IN3 n2531 n121 n260 n97 n470 VDD VSS OAI221_X1 
XU49 IN3 n2531 n122 n259 n98 n471 VDD VSS OAI221_X1 
XU48 IN3 n2531 n118 n260 n94 n467 VDD VSS OAI221_X1 
XU47 IN3 n2531 n94 n260 n65 n443 VDD VSS OAI221_X1 
XU46 IN3 n2531 n597 n259 n90 n463 VDD VSS OAI221_X1 
XU45 IN3 n2531 n115 n259 n91 n464 VDD VSS OAI221_X1 
XU44 IN3 n2531 n110 n260 n86 n459 VDD VSS OAI221_X1 
XU43 IN3 n2531 n609 n259 n1300 n465 VDD VSS OAI221_X1 
XU42 IN3 n2531 n111 n259 n87 n460 VDD VSS OAI221_X1 
XU41 IN3 n2531 n117 n259 n93 n466 VDD VSS OAI221_X1 
XU40 IN3 n2531 n112 n259 n88 n461 VDD VSS OAI221_X1 
XU39 IN3 n2531 n113 n259 n89 n462 VDD VSS OAI221_X1 
XU38 IN2 n255 n140 n258 n124 n376 VDD VSS OAI221_X1 
XU37 n252 n1080 N2610 VDD VSS NOR2_X1 
XU36 n252 n331 N2600 VDD VSS NOR2_X1 
XU35 n252 n333 N2590 VDD VSS NOR2_X1 
XU34 n252 n1090 N2580 VDD VSS NOR2_X1 
XU33 n252 n1095 N2570 VDD VSS NOR2_X1 
XU32 n252 n1100 N2560 VDD VSS NOR2_X1 
XU31 n252 n1105 N2550 VDD VSS NOR2_X1 
XU19 IN0 n255 n188 VDD VSS NAND2_X1 
XU18 n188 n258 VDD VSS BUF_X2 
XU17 n187 n257 VDD VSS BUF_X2 
XU15 n187 n255 VDD VSS BUF_X2 
XU14 n187 n254 VDD VSS BUF_X2 
XU13 n187 n2531 VDD VSS BUF_X2 
XU441 n373 n374 n372 VDD VSS XOR2_X1 
XU440 n369 n370 n368 VDD VSS XOR2_X1 
XU439 n365 n366 n364 VDD VSS XOR2_X1 
XU438 n361 n362 n360 VDD VSS XOR2_X1 
XU437 n357 n358 n356 VDD VSS XOR2_X1 
XU436 n353 n354 n352 VDD VSS XOR2_X1 
XU435 n83 z1[45] n220 VDD VSS XOR2_X1 
XU434 n201 n220 n351 VDD VSS XOR2_X1 
XU433 n350 n351 n349 VDD VSS XOR2_X1 
XU432 n81 z1[46] n219 VDD VSS XOR2_X1 
XU431 n200 n219 n348 VDD VSS XOR2_X1 
XU430 n347 n348 n346 VDD VSS XOR2_X1 
XU429 n79 z1[47] n218 VDD VSS XOR2_X1 
XU428 n199 n218 n345 VDD VSS XOR2_X1 
XU427 n344 n345 n343 VDD VSS XOR2_X1 
XU426 n77 z1[48] n217 VDD VSS XOR2_X1 
XU425 n198 n217 n342 VDD VSS XOR2_X1 
XU424 n232 n342 n341 VDD VSS XOR2_X1 
XU423 n75 z1[49] n216 VDD VSS XOR2_X1 
XU169 IN2 n255 n161 n258 n1573 n397 VDD VSS OAI221_X1 
XU168 IN2 n255 n1573 n258 n135 n384 VDD VSS OAI221_X1 
XU167 IN2 n255 n167 n258 n154 n403 VDD VSS OAI221_X1 
XU166 IN2 n255 n141 n258 n126 n377 VDD VSS OAI221_X1 
XU165 IN2 n255 n173 n258 n160 n409 VDD VSS OAI221_X1 
XU164 IN2 n255 n160 n258 n147 n396 VDD VSS OAI221_X1 
XU163 IN2 n255 n147 n258 n134 n383 VDD VSS OAI221_X1 
XU162 IN0 n255 n166 n260 n153 n402 VDD VSS OAI221_X1 
XU161 IN2 n255 n153 n140 n258 n389 VDD VSS OAI221_X1 
XU160 IN0 n255 n172 n260 n774 n408 VDD VSS OAI221_X1 
XU159 IN0 n255 n774 n260 n146 n395 VDD VSS OAI221_X1 
XU158 IN0 n257 n146 n261 n133 n382 VDD VSS OAI221_X1 
XU157 IN0 n257 n165 n261 n152 n401 VDD VSS OAI221_X1 
XU156 IN0 n257 n152 n261 n139 n388 VDD VSS OAI221_X1 
XU155 n225 n623 VDD VSS INV_X1 
XU154 IN3 n623 n2531 n259 n735 n496 VDD VSS OAI221_X1 
XU153 IN2 n231 n255 n258 n698 n550 VDD VSS OAI221_X1 
XU152 IN2 n226 n255 n258 n719 n545 VDD VSS OAI221_X1 
XU151 IN0 n229 n254 n261 n1886 n548 VDD VSS OAI221_X1 
XU150 n221 n619 VDD VSS INV_X1 
XU149 IN2 n619 n255 n260 n119 n492 VDD VSS OAI221_X1 
XU148 n224 n622 VDD VSS INV_X1 
XU147 IN3 n622 n2531 n259 n122 n495 VDD VSS OAI221_X1 
XU146 IN3 n206 n2531 n259 n104 n477 VDD VSS OAI221_X1 
XU145 IN2 n202 n255 n260 n100 n473 VDD VSS OAI221_X1 
XU144 IN3 n203 n2531 n259 n101 n474 VDD VSS OAI221_X1 
XU143 IN3 n218 n2531 n259 n609 n489 VDD VSS OAI221_X1 
XU142 IN3 n204 n2531 n259 n102 n475 VDD VSS OAI221_X1 
XU141 IN0 n200 n257 n259 n183 n432 VDD VSS OAI221_X1 
XU140 rstn n198 n254 n258 n667 n430 VDD VSS OAI221_X1 
XU139 IN2 n197 n255 n258 n1581 n429 VDD VSS OAI221_X1 
XU138 n261 n27 n254 n34 n523 VDD VSS OAI22_X1 
XU137 n261 n30 n254 n37 n526 VDD VSS OAI22_X1 
XU136 n261 n23 n254 n30 n519 VDD VSS OAI22_X1 
XU135 n261 n700 n254 n40 n529 VDD VSS OAI22_X1 
XU134 n261 n701 n254 n700 n522 VDD VSS OAI22_X1 
XU133 n261 n29 n254 n36 n525 VDD VSS OAI22_X1 
XU132 n260 n32 n257 n39 n528 VDD VSS OAI22_X1 
XU131 n260 n25 n2531 n32 n521 VDD VSS OAI22_X1 
XU130 n260 n18 n2531 n25 n514 VDD VSS OAI22_X1 
XU129 n260 n28 n255 n35 n524 VDD VSS OAI22_X1 
XU128 n258 n21 n254 n28 n517 VDD VSS OAI22_X1 
XU127 n261 n729 n254 n727 n527 VDD VSS OAI22_X1 
XU126 n260 n70 n2531 n99 n448 VDD VSS OAI22_X1 
XU125 n260 n56 n2531 n85 n434 VDD VSS OAI22_X1 
XU124 n260 n66 n255 n95 n444 VDD VSS OAI22_X1 
XU123 n260 n77 n255 n105 n454 VDD VSS OAI22_X1 
XU122 n259 n79 n2531 n2001 n455 VDD VSS OAI22_X1 
XU121 n259 n68 n2531 n97 n446 VDD VSS OAI22_X1 
XU120 n259 n81 n257 n107 n456 VDD VSS OAI22_X1 
XU119 n259 n69 n257 n98 n447 VDD VSS OAI22_X1 
XU118 n259 n83 n257 n108 n457 VDD VSS OAI22_X1 
XU117 n260 n75 n2531 n104 n453 VDD VSS OAI22_X1 
XU116 n260 n71 n255 n100 n449 VDD VSS OAI22_X1 
XU115 n259 n62 n2531 n91 n440 VDD VSS OAI22_X1 
XU114 n259 n72 n2531 n101 n450 VDD VSS OAI22_X1 
XU113 n259 n58 n2531 n87 n436 VDD VSS OAI22_X1 
XU112 n259 n73 n2531 n102 n451 VDD VSS OAI22_X1 
XU111 n259 n59 n257 n88 n437 VDD VSS OAI22_X1 
XU110 n259 n74 n257 n103 n452 VDD VSS OAI22_X1 
XU109 n259 n60 n2531 n89 n438 VDD VSS OAI22_X1 
XU108 n259 n1396 n257 n184 n420 VDD VSS OAI22_X1 
XU107 n260 n1152 n257 n1418 n413 VDD VSS OAI22_X1 
XU106 n259 n170 n257 n183 n419 VDD VSS OAI22_X1 
XU105 n259 n1491 n257 n182 n418 VDD VSS OAI22_X1 
XU104 n258 n1537 n254 n667 n417 VDD VSS OAI22_X1 
XU103 n258 n161 n255 n174 n410 VDD VSS OAI22_X1 
XU102 n258 n167 n255 n1581 n416 VDD VSS OAI22_X1 
XU101 n258 n166 n254 n179 n415 VDD VSS OAI22_X1 
XU100 n259 n165 n257 n178 n414 VDD VSS OAI22_X1 
XU99 n258 n1646 n255 n1640 n544 VDD VSS OAI22_X1 
XU98 n258 n34 n254 n41 n530 VDD VSS OAI22_X1 
XU97 n261 n37 n254 n44 n533 VDD VSS OAI22_X1 
XU96 n258 n40 n255 n47 n536 VDD VSS OAI22_X1 
XU95 n261 n36 n254 n43 n532 VDD VSS OAI22_X1 
XU94 n260 n39 n257 n46 n535 VDD VSS OAI22_X1 
XU93 n260 n11 n257 n18 n507 VDD VSS OAI22_X1 
XU92 n258 n35 n255 n42 n531 VDD VSS OAI22_X1 
XU91 n261 n727 n257 n726 n534 VDD VSS OAI22_X1 
XU90 n261 n144 n257 n157 n393 VDD VSS OAI22_X1 
XU89 n258 n142 n254 n155 n391 VDD VSS OAI22_X1 
XU88 n258 n141 n255 n154 n390 VDD VSS OAI22_X1 
XU87 n222 n620 VDD VSS INV_X1 
XU86 IN2 n620 n255 n260 n120 n493 VDD VSS OAI221_X1 
XU85 n223 n621 VDD VSS INV_X1 
XU84 IN3 n621 n2531 n260 n121 n494 VDD VSS OAI221_X1 
XU83 IN3 n220 n2531 n260 n118 n491 VDD VSS OAI221_X1 
XU82 IN3 n216 n2531 n259 n597 n487 VDD VSS OAI221_X1 
XU81 IN3 n219 n2531 n259 n117 n490 VDD VSS OAI221_X1 
XU80 IN3 n205 n257 n259 n103 n476 VDD VSS OAI221_X1 
XU79 IN0 n254 n27 n261 n20 n516 VDD VSS OAI221_X1 
XU78 IN0 n254 n51 n261 n44 n540 VDD VSS OAI221_X1 
XU77 IN0 n254 n701 n261 n703 n515 VDD VSS OAI221_X1 
XU262 z2_next[20] z3_next[20] n320 VDD VSS XNOR2_X1 
XU261 n320 n206 n319 VDD VSS XNOR2_X1 
XU260 n185 n1053 N266 VDD VSS NOR2_X1 
XU259 z2_next[19] z3_next[19] n322 VDD VSS XNOR2_X1 
XU258 n322 n207 n321 VDD VSS XNOR2_X1 
XU257 n185 n1058 N265 VDD VSS NOR2_X1 
XU256 z3_next[18] n189 n324 VDD VSS XNOR2_X1 
XU255 n324 n208 n323 VDD VSS XNOR2_X1 
XU254 n185 n1063 N264 VDD VSS NOR2_X1 
XU253 z3_next[17] n190 n326 VDD VSS XNOR2_X1 
XU252 n326 n209 n325 VDD VSS XNOR2_X1 
XU251 n252 n1068 N263 VDD VSS NOR2_X1 
XU250 z3_next[16] n191 n328 VDD VSS XNOR2_X1 
XU249 n328 n210 n327 VDD VSS XNOR2_X1 
XU248 n252 n1073 N262 VDD VSS NOR2_X1 
XU247 z3_next[39] z3_next[63] n344 VDD VSS XNOR2_X1 
XU246 n252 n1110 N2540 VDD VSS NOR2_X1 
XU245 z3_next[38] z3_next[62] n347 VDD VSS XNOR2_X1 
XU244 n252 n1115 N253 VDD VSS NOR2_X1 
XU243 z3_next[37] z3_next[61] n350 VDD VSS XNOR2_X1 
XU242 n252 n1120 N2520 VDD VSS NOR2_X1 
XU241 n140 n355 n354 VDD VSS XNOR2_X1 
XU240 z2_next[44] n221 n353 VDD VSS XNOR2_X1 
XU239 n252 n1124 N251 VDD VSS NOR2_X1 
XU238 n141 n359 n358 VDD VSS XNOR2_X1 
XU237 z2_next[43] n222 n357 VDD VSS XNOR2_X1 
XU236 n252 n1129 N2500 VDD VSS NOR2_X1 
XU235 z2_next[42] n223 n361 VDD VSS XNOR2_X1 
XU234 n142 n363 n362 VDD VSS XNOR2_X1 
XU233 n252 n1134 N249 VDD VSS NOR2_X1 
XU232 n143 n367 n366 VDD VSS XNOR2_X1 
XU231 z2_next[41] n224 n365 VDD VSS XNOR2_X1 
XU230 n250 n1139 N2480 VDD VSS NOR2_X1 
XU229 n144 n371 n370 VDD VSS XNOR2_X1 
XU228 z2_next[40] n225 n369 VDD VSS XNOR2_X1 
XU227 n246 n1144 N247 VDD VSS NOR2_X1 
XU226 n1152 n375 n374 VDD VSS XNOR2_X1 
XU225 n576 n244 n373 VDD VSS XNOR2_X1 
XU224 n185 n1148 N2460 VDD VSS NOR2_X1 
XU222 n261 n732 n254 n24 n513 VDD VSS OAI22_X1 
XU221 n261 n16 n254 n23 n512 VDD VSS OAI22_X1 
XU220 n261 n14 n254 n21 n510 VDD VSS OAI22_X1 
XU219 ce IN3 n187 VDD VSS NAND2_X1 
XU218 n258 n1640 n232 n255 n551 VDD VSS OAI22_X1 
XU217 n261 n1681 n228 n254 n547 VDD VSS OAI22_X1 
XU216 n261 n1765 n227 n254 n546 VDD VSS OAI22_X1 
XU215 n260 n53 n230 n255 n549 VDD VSS OAI22_X1 
XU214 n259 n2001 n208 n2531 n479 VDD VSS OAI22_X1 
XU213 n259 n107 n209 n2531 n480 VDD VSS OAI22_X1 
XU212 n259 n587 n210 n257 n481 VDD VSS OAI22_X1 
XU211 n259 n115 n217 n2531 n488 VDD VSS OAI22_X1 
XU210 n260 n110 n212 n2531 n483 VDD VSS OAI22_X1 
XU209 n261 n1418 n194 n257 n426 VDD VSS OAI22_X1 
XU208 n261 n176 n193 n257 n425 VDD VSS OAI22_X1 
XU207 n191 n624 VDD VSS INV_X1 
XU206 n258 n174 n624 n255 n423 VDD VSS OAI22_X1 
XU205 n260 n109 n211 n2531 n482 VDD VSS OAI22_X1 
XU204 n260 n105 n207 n255 n478 VDD VSS OAI22_X1 
XU203 n259 n111 n213 n2531 n484 VDD VSS OAI22_X1 
XU202 n259 n112 n214 n2531 n485 VDD VSS OAI22_X1 
XU201 n259 n113 n215 n257 n486 VDD VSS OAI22_X1 
XU200 n259 n184 n201 n257 n433 VDD VSS OAI22_X1 
XU199 n259 n182 n199 n257 n431 VDD VSS OAI22_X1 
XU198 n258 n175 n192 n254 n424 VDD VSS OAI22_X1 
XU197 n190 n625 VDD VSS INV_X1 
XU196 n258 n173 n625 n255 n422 VDD VSS OAI22_X1 
XU195 n258 n179 n196 n254 n428 VDD VSS OAI22_X1 
XU194 n189 n626 VDD VSS INV_X1 
XU193 n260 n172 n626 n255 n421 VDD VSS OAI22_X1 
XU192 n261 n178 n195 n257 n427 VDD VSS OAI22_X1 
XU191 IN3 n2531 n90 n260 n1974 n439 VDD VSS OAI221_X1 
XU190 IN3 n2531 n86 n260 n57 n435 VDD VSS OAI221_X1 
XU189 IN3 n2531 n1300 n259 n63 n441 VDD VSS OAI221_X1 
XU188 IN3 n2531 n93 n259 n64 n442 VDD VSS OAI221_X1 
XU187 IN3 n257 n1396 n259 n643 n407 VDD VSS OAI221_X1 
XU186 IN0 n257 n643 n259 n1406 n394 VDD VSS OAI221_X1 
XU185 IN0 n257 n1406 n261 n132 n381 VDD VSS OAI221_X1 
XU184 IN0 n257 n1152 n261 n151 n400 VDD VSS OAI221_X1 
XU183 IN0 n257 n151 n261 n138 n387 VDD VSS OAI221_X1 
XU182 IN3 n257 n170 n259 n157 n406 VDD VSS OAI221_X1 
XU181 IN0 n257 n144 n261 n131 n380 VDD VSS OAI221_X1 
XU180 IN0 n257 n176 n259 n1470 n412 VDD VSS OAI221_X1 
XU179 IN0 n257 n1470 n259 n150 n399 VDD VSS OAI221_X1 
XU178 IN0 n257 n150 n261 n137 n386 VDD VSS OAI221_X1 
XU177 IN3 n257 n1491 n259 n156 n405 VDD VSS OAI221_X1 
XU176 IN0 n257 n156 n261 n143 n392 VDD VSS OAI221_X1 
XU175 IN0 n254 n143 n261 n130 n379 VDD VSS OAI221_X1 
XU174 rstn n254 n175 n258 n162 n411 VDD VSS OAI221_X1 
XU173 rstn n254 n162 n258 n149 n398 VDD VSS OAI221_X1 
XU172 rstn n254 n149 n258 n136 n385 VDD VSS OAI221_X1 
XU171 rstn n254 n1537 n258 n155 n404 VDD VSS OAI221_X1 
XU170 rstn n254 n142 n258 n128 n378 VDD VSS OAI221_X1 
XU355 n20 z2_next[51] n25800 VDD VSS XNOR2_X1 
XU354 z1_next[51] n25800 n25700 VDD VSS XNOR2_X1 
XU353 n185 n878 N297 VDD VSS NOR2_X1 
XU352 n21 z2_next[50] n26000 VDD VSS XNOR2_X1 
XU351 z1_next[50] n26000 n25900 VDD VSS XNOR2_X1 
XU350 n252 n886 N296 VDD VSS NOR2_X1 
XU349 n22 z2_next[49] n2620 VDD VSS XNOR2_X1 
XU348 z1_next[49] n2620 n26100 VDD VSS XNOR2_X1 
XU347 n185 n890 N295 VDD VSS NOR2_X1 
XU346 n23 z2_next[48] n2640 VDD VSS XNOR2_X1 
XU345 z1_next[48] n2640 n2630 VDD VSS XNOR2_X1 
XU344 n185 n896 N294 VDD VSS NOR2_X1 
XU343 n24 z2_next[47] n2660 VDD VSS XNOR2_X1 
XU342 z1_next[47] n2660 n2650 VDD VSS XNOR2_X1 
XU341 n248 n902 N293 VDD VSS NOR2_X1 
XU340 n25 z2_next[46] n2680 VDD VSS XNOR2_X1 
XU339 z1_next[46] n2680 n2670 VDD VSS XNOR2_X1 
XU338 n248 n908 N292 VDD VSS NOR2_X1 
XU337 n26 z2_next[45] n2700 VDD VSS XNOR2_X1 
XU336 z1_next[45] n2700 n2690 VDD VSS XNOR2_X1 
XU335 n246 n914 N291 VDD VSS NOR2_X1 
XU334 n27 z2_next[44] n2720 VDD VSS XNOR2_X1 
XU333 z1_next[44] n2720 n2710 VDD VSS XNOR2_X1 
XU332 n246 n920 N290 VDD VSS NOR2_X1 
XU331 n28 z2_next[43] n2740 VDD VSS XNOR2_X1 
XU330 z1_next[43] n2740 n2730 VDD VSS XNOR2_X1 
XU329 n246 n926 N289 VDD VSS NOR2_X1 
XU328 n29 z2_next[42] n2760 VDD VSS XNOR2_X1 
XU327 z1_next[42] n2760 n2750 VDD VSS XNOR2_X1 
XU326 n246 n932 N288 VDD VSS NOR2_X1 
XU325 n30 z2_next[41] n2780 VDD VSS XNOR2_X1 
XU324 z1_next[41] n2780 n2770 VDD VSS XNOR2_X1 
XU323 n246 n938 N287 VDD VSS NOR2_X1 
XU322 n31 z2_next[40] n2800 VDD VSS XNOR2_X1 
XU321 z1_next[40] n2800 n2790 VDD VSS XNOR2_X1 
XU320 n246 n940 N286 VDD VSS NOR2_X1 
XU319 n32 z2_next[39] n2820 VDD VSS XNOR2_X1 
XU318 z1_next[39] n2820 n2810 VDD VSS XNOR2_X1 
XU317 n246 n946 N285 VDD VSS NOR2_X1 
XU316 n33 z2_next[38] n2840 VDD VSS XNOR2_X1 
XU315 z1_next[38] n2840 n2830 VDD VSS XNOR2_X1 
XU314 n246 n952 N284 VDD VSS NOR2_X1 
XU313 n34 z2_next[37] n2860 VDD VSS XNOR2_X1 
XU312 z1_next[37] n2860 n2850 VDD VSS XNOR2_X1 
XU311 n246 n958 N283 VDD VSS NOR2_X1 
XU310 n35 z2_next[36] n2880 VDD VSS XNOR2_X1 
XU309 z1_next[36] n2880 n2870 VDD VSS XNOR2_X1 
XU308 n246 n964 N282 VDD VSS NOR2_X1 
XU307 n36 z2_next[35] n2900 VDD VSS XNOR2_X1 
XU306 z1_next[35] n2900 n2890 VDD VSS XNOR2_X1 
XU305 n246 n970 N281 VDD VSS NOR2_X1 
XU304 n37 z2_next[34] n2920 VDD VSS XNOR2_X1 
XU303 z1_next[34] n2920 n2910 VDD VSS XNOR2_X1 
XU302 n246 n977 N280 VDD VSS NOR2_X1 
XU301 n38 z2_next[33] n2940 VDD VSS XNOR2_X1 
XU300 z1_next[33] n2940 n2930 VDD VSS XNOR2_X1 
XU299 n246 n981 N279 VDD VSS NOR2_X1 
XU298 n39 z2_next[32] n2960 VDD VSS XNOR2_X1 
XU297 z1_next[32] n2960 n2950 VDD VSS XNOR2_X1 
XU296 n246 n987 N278 VDD VSS NOR2_X1 
XU295 n40 z2_next[31] n2980 VDD VSS XNOR2_X1 
XU294 z1_next[31] n2980 n2970 VDD VSS XNOR2_X1 
XU293 n185 n993 N277 VDD VSS NOR2_X1 
XU292 n41 z2_next[30] n3000 VDD VSS XNOR2_X1 
XU291 z1_next[30] n3000 n2990 VDD VSS XNOR2_X1 
XU290 n185 n999 N276 VDD VSS NOR2_X1 
XU289 n42 z2_next[29] n3020 VDD VSS XNOR2_X1 
XU288 z1_next[29] n3020 n3010 VDD VSS XNOR2_X1 
XU287 n185 n1007 N275 VDD VSS NOR2_X1 
XU286 n43 z2_next[28] n3040 VDD VSS XNOR2_X1 
XU285 z1_next[28] n3040 n3030 VDD VSS XNOR2_X1 
XU284 n185 n1011 N274 VDD VSS NOR2_X1 
XU283 n44 z2_next[27] n3060 VDD VSS XNOR2_X1 
XU282 z1_next[27] n3060 n3050 VDD VSS XNOR2_X1 
XU281 n185 n1016 N273 VDD VSS NOR2_X1 
XU280 n45 z2_next[26] n3080 VDD VSS XNOR2_X1 
XU279 z1_next[26] n3080 n3070 VDD VSS XNOR2_X1 
XU278 n185 n1020 N272 VDD VSS NOR2_X1 
XU277 n46 z2_next[25] n310 VDD VSS XNOR2_X1 
XU276 z1_next[25] n310 n3090 VDD VSS XNOR2_X1 
XU275 n185 n1025 N271 VDD VSS NOR2_X1 
XU274 z2_next[24] z3_next[24] n312 VDD VSS XNOR2_X1 
XU273 n312 n202 n311 VDD VSS XNOR2_X1 
XU272 n185 n1031 N270 VDD VSS NOR2_X1 
XU271 z2_next[23] z3_next[23] n314 VDD VSS XNOR2_X1 
XU270 n314 n203 n313 VDD VSS XNOR2_X1 
XU269 n185 n1037 N269 VDD VSS NOR2_X1 
XU268 z2_next[22] z3_next[22] n316 VDD VSS XNOR2_X1 
XU267 n316 n204 n315 VDD VSS XNOR2_X1 
XU266 n185 n1042 N268 VDD VSS NOR2_X1 
XU265 z2_next[21] z3_next[21] n318 VDD VSS XNOR2_X1 
XU264 n318 n205 n317 VDD VSS XNOR2_X1 
XU263 n185 n1047 N267 VDD VSS NOR2_X1 
XU467 n13 z3_next[34] n363 VDD VSS XNOR2_X1 
XU466 n12 z3_next[35] n359 VDD VSS XNOR2_X1 
XU465 n1797 z3_next[32] n371 VDD VSS XNOR2_X1 
XU464 n11 z3_next[36] n355 VDD VSS XNOR2_X1 
XU463 n14 z3_next[33] n367 VDD VSS XNOR2_X1 
XU462 n16 z3_next[31] n375 VDD VSS XNOR2_X1 
XU461 z3[62] z3_next[45] n227 VDD VSS XNOR2_X1 
XU460 z3[61] z3_next[44] n228 VDD VSS XNOR2_X1 
XU459 z3[59] z3_next[42] n230 VDD VSS XNOR2_X1 
XU458 z3[57] z3_next[40] n232 VDD VSS XNOR2_X1 
XU457 n130 n149 n192 VDD VSS XNOR2_X1 
XU456 n131 n150 n193 VDD VSS XNOR2_X1 
XU455 n132 n151 n194 VDD VSS XNOR2_X1 
XU454 n133 n152 n195 VDD VSS XNOR2_X1 
XU453 n134 n153 n196 VDD VSS XNOR2_X1 
XU452 n137 n156 n199 VDD VSS XNOR2_X1 
XU451 n139 n158 n201 VDD VSS XNOR2_X1 
XU450 z3[63] z3_next[46] n226 VDD VSS XNOR2_X1 
XU449 z3[60] z3_next[43] n229 VDD VSS XNOR2_X1 
XU448 z3[58] z3_next[41] n231 VDD VSS XNOR2_X1 
XU447 n135 n154 n197 VDD VSS XNOR2_X1 
XU446 n136 n155 n198 VDD VSS XNOR2_X1 
XU445 n138 n157 n200 VDD VSS XNOR2_X1 
XU444 n66 n1974 n207 VDD VSS XNOR2_X1 
XU443 n68 n63 n209 VDD VSS XNOR2_X1 
XU442 n69 n64 n210 VDD VSS XNOR2_X1 
XU405 n67 n62 n208 VDD VSS XNOR2_X1 
XU404 z2[63] n146 n189 VDD VSS XNOR2_X1 
XU403 z2[62] n147 n190 VDD VSS XNOR2_X1 
XU402 z2[61] n1573 n191 VDD VSS XNOR2_X1 
XU401 z1[43] n86 n222 VDD VSS XNOR2_X1 
XU400 z1[44] n85 n221 VDD VSS XNOR2_X1 
XU399 z1[42] n87 n223 VDD VSS XNOR2_X1 
XU398 z1[41] n88 n224 VDD VSS XNOR2_X1 
XU397 z1[40] n89 n225 VDD VSS XNOR2_X1 
XU396 n65 n60 n206 VDD VSS XNOR2_X1 
XU395 n1974 n56 n202 VDD VSS XNOR2_X1 
XU394 n63 n58 n204 VDD VSS XNOR2_X1 
XU393 n64 n59 n205 VDD VSS XNOR2_X1 
XU392 n62 n57 n203 VDD VSS XNOR2_X1 
XU391 n90 z2_next[58] n244 VDD VSS XNOR2_X1 
XU390 n806 z2_next[63] n234 VDD VSS XNOR2_X1 
XU389 n576 n234 n233 VDD VSS XNOR2_X1 
XU388 n252 n808 N3091 VDD VSS NOR2_X1 
XU387 n9 z2_next[62] n236 VDD VSS XNOR2_X1 
XU386 z1_next[62] n236 n235 VDD VSS XNOR2_X1 
XU385 n252 n814 N3081 VDD VSS NOR2_X1 
XU384 n10 z2_next[61] n238 VDD VSS XNOR2_X1 
XU383 z1_next[61] n238 n237 VDD VSS XNOR2_X1 
XU382 n252 n820 N3071 VDD VSS NOR2_X1 
XU381 n11 z2_next[60] n240 VDD VSS XNOR2_X1 
XU380 z1_next[60] n240 n239 VDD VSS XNOR2_X1 
XU379 n252 n826 N3061 VDD VSS NOR2_X1 
XU378 n12 z2_next[59] n242 VDD VSS XNOR2_X1 
XU377 z1_next[59] n242 n241 VDD VSS XNOR2_X1 
XU376 n252 n832 N3051 VDD VSS NOR2_X1 
XU375 z3_next[58] n244 n243 VDD VSS XNOR2_X1 
XU374 n252 n838 N3041 VDD VSS NOR2_X1 
XU373 n14 z2_next[57] n24600 VDD VSS XNOR2_X1 
XU372 z1_next[57] n24600 n245 VDD VSS XNOR2_X1 
XU371 n185 n843 N303 VDD VSS NOR2_X1 
XU370 n1797 z2_next[56] n24800 VDD VSS XNOR2_X1 
XU369 z1_next[56] n24800 n2470 VDD VSS XNOR2_X1 
XU368 n185 n848 N302 VDD VSS NOR2_X1 
XU367 n16 z2_next[55] n25000 VDD VSS XNOR2_X1 
XU366 z1_next[55] n25000 n2490 VDD VSS XNOR2_X1 
XU365 n185 n854 N301 VDD VSS NOR2_X1 
XU364 n17 z2_next[54] n25200 VDD VSS XNOR2_X1 
XU363 z1_next[54] n25200 n2510 VDD VSS XNOR2_X1 
XU362 n185 n860 N300 VDD VSS NOR2_X1 
XU361 n18 z2_next[53] n25400 VDD VSS XNOR2_X1 
XU360 z1_next[53] n25400 n2530 VDD VSS XNOR2_X1 
XU359 n185 n868 N299 VDD VSS NOR2_X1 
XU358 n19 z2_next[52] n25600 VDD VSS XNOR2_X1 
XU357 z1_next[52] n25600 n25500 VDD VSS XNOR2_X1 
XU356 n185 n874 N298 VDD VSS NOR2_X1 
XCLKBUF_X1_G2B1I1 n78 n78_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I2 n78 n78_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I4 n78 n78_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I5 n78 n78_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I6 n78 n78_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I7 n78 n78_G2B1I7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I8 n78 n78_G2B1I8 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I11 n125 n125_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I31 n125 n125_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I41 n125 n125_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I51 n125 n125_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I61 n125 n125_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I22 n84 n84_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I32 n84 n84_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I42 n84 n84_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I52 n84 n84_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I62 n84 n84_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I13 n76 n76_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I33 n76 n76_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I43 n76 n76_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I24 clk_G1B1I2 n82_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I34 clk_G1B1I2 n82_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I44 clk_G1B1I2 n82_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I53 clk_G1B1I2 n82_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I63 clk_G1B1I2 n82_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I71 clk_G1B1I2 n82_G2B1I7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I81 clk_G1B1I2 n82_G2B1I8 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I15 n80 n80_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I25 n80 n80_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I45 n80 n80_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I54 n80 n80_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I64 n80 n80_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I72 n80 n80_G2B1I7 VDD VSS CLKBUF_X1 
XU6 clk_cts_3 n125 VDD VSS CLKBUF_X1 
XCLKBUF_X3_G1B1I6 clk clk_G1B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X3_G1B1I3 clk clk_G1B1I3 VDD VSS CLKBUF_X1 
XU1 clk_G1B1I3 n76 VDD VSS CLKBUF_X1 
XCLKBUF_X2_G1B1I2 clk clk_G1B1I2 VDD VSS CLKBUF_X1 
XU5 clk_G1B1I3 n84 VDD VSS CLKBUF_X1 
XU2 clk_G1B1I6 n78 VDD VSS CLKBUF_X1 
XU3 clk_G1B1I6 n80 VDD VSS CLKBUF_X1 
XU4 n810 n304 VDD VSS BUF_X1 
XU8 n841 n305 VDD VSS BUF_X1 
XU23 n876 n306 VDD VSS BUF_X1 
XU24 n572 n307 VDD VSS BUF_X1 
XU25 n991 n308 VDD VSS BUF_X1 
XU26 n574 n309 VDD VSS BUF_X1 
XU27 n1018 n552 VDD VSS BUF_X1 
XU28 n1107 n553 VDD VSS BUF_X1 
XU29 n575 n554 VDD VSS BUF_X1 
XU30 n1150 n555 VDD VSS BUF_X1 
XU223 n1901 n556 VDD VSS BUF_X1 
XU468 n61 n1973 VDD VSS INV_X16 
XU469 n148 n1572 VDD VSS INV_X16 
XU470 n343 n1108 VDD VSS BUF_X1 
XU471 n3050 n1012 VDD VSS BUF_X1 
XU472 n990 n991 VDD VSS INV_X8 
XU473 n961 n962 VDD VSS INV_X8 
XU474 n911 n912 VDD VSS INV_X2 
XU475 n753 n557 VDD VSS INV_X1 
XU476 n557 n558 VDD VSS INV_X8 
XU477 n758 n559 VDD VSS BUF_X1 
XU478 n763 n560 VDD VSS CLKBUF_X1 
XU479 n773 n561 VDD VSS BUF_X1 
XU480 n772 n562 VDD VSS CLKBUF_X1 
XU481 n779 n563 VDD VSS BUF_X1 
XU482 n784 n564 VDD VSS BUF_X1 
XU483 n789 n565 VDD VSS BUF_X1 
XU484 n786 n566 VDD VSS CLKBUF_X1 
XU485 n794 n567 VDD VSS BUF_X1 
XU486 n791 n568 VDD VSS CLKBUF_X1 
XU487 n799 n569 VDD VSS INV_X1 
XU488 n569 n570 VDD VSS INV_X32 
XU489 n804 n571 VDD VSS BUF_X1 
XU490 n912 n572 VDD VSS BUF_X1 
XU491 n930 n573 VDD VSS BUF_X1 
XU492 n1014 n574 VDD VSS BUF_X1 
XU493 n1112 n575 VDD VSS BUF_X1 
XU494 z1_next[63] n576 VDD VSS CLKBUF_X1 
XU495 n1157 n577 VDD VSS BUF_X1 
XU496 n1162 n578 VDD VSS BUF_X1 
XU497 n1159 n579 VDD VSS CLKBUF_X1 
XU498 n1167 n580 VDD VSS INV_X1 
XU499 n580 n581 VDD VSS INV_X8 
XU500 n1178 n582 VDD VSS BUF_X1 
XU501 n1183 n583 VDD VSS BUF_X1 
XU502 n1188 n584 VDD VSS BUF_X1 
XU503 n1186 n585 VDD VSS CLKBUF_X1 
XU504 n1193 n586 VDD VSS BUF_X1 
XU505 n108 n587 VDD VSS CLKBUF_X1 
XU506 n1198 n588 VDD VSS CLKBUF_X1 
XU507 n1203 n589 VDD VSS BUF_X1 
XU508 n1208 n590 VDD VSS BUF_X1 
XU509 n1213 n591 VDD VSS BUF_X1 
XU510 n1218 n592 VDD VSS INV_X1 
XU511 n592 n593 VDD VSS INV_X8 
XU512 n1223 n594 VDD VSS BUF_X1 
XU513 n1220 n595 VDD VSS CLKBUF_X1 
XU514 n1233 n596 VDD VSS BUF_X1 
XU515 n114 n597 VDD VSS CLKBUF_X1 
XU516 n1243 n598 VDD VSS BUF_X1 
XU517 n1248 n599 VDD VSS BUF_X1 
XU518 n1246 n600 VDD VSS CLKBUF_X1 
XU519 n1259 n601 VDD VSS BUF_X1 
XU520 n1270 n602 VDD VSS BUF_X1 
XU521 n1268 n603 VDD VSS CLKBUF_X1 
XU522 n1275 n604 VDD VSS BUF_X1 
XU523 n1280 n605 VDD VSS BUF_X1 
XU524 n1285 n606 VDD VSS BUF_X1 
XU525 n1290 n607 VDD VSS CLKBUF_X1 
XU526 n1299 n608 VDD VSS BUF_X1 
XU527 n116 n609 VDD VSS CLKBUF_X1 
XU528 n1298 n610 VDD VSS CLKBUF_X1 
XU529 n1305 n611 VDD VSS BUF_X1 
XU530 n1310 n612 VDD VSS INV_X1 
XU531 n612 n613 VDD VSS INV_X8 
XU532 n1315 n614 VDD VSS BUF_X1 
XU533 n1320 n615 VDD VSS CLKBUF_X1 
XU534 n1325 n616 VDD VSS BUF_X1 
XU535 n1330 n617 VDD VSS BUF_X1 
XU536 n1328 n618 VDD VSS CLKBUF_X1 
XU537 n1335 n627 VDD VSS BUF_X1 
XU538 n1340 n628 VDD VSS BUF_X1 
XU539 n1345 n629 VDD VSS BUF_X1 
XU540 n1350 n630 VDD VSS BUF_X1 
XU541 n1347 n631 VDD VSS CLKBUF_X1 
XU542 n1355 n632 VDD VSS BUF_X1 
XU543 n1360 n633 VDD VSS CLKBUF_X1 
XU544 n1365 n634 VDD VSS BUF_X1 
XU545 n1370 n635 VDD VSS CLKBUF_X1 
XU546 n1373 n636 VDD VSS BUF_X1 
XU547 n1375 n637 VDD VSS CLKBUF_X1 
XU548 n1380 n638 VDD VSS BUF_X1 
XU549 n1385 n639 VDD VSS BUF_X1 
XU550 n1395 n640 VDD VSS INV_X1 
XU551 n640 n641 VDD VSS INV_X32 
XU552 n1405 n642 VDD VSS BUF_X1 
XU553 n158 n643 VDD VSS BUF_X1 
XU554 n1404 n644 VDD VSS CLKBUF_X1 
XU555 n1411 n645 VDD VSS BUF_X1 
XU556 n1427 n646 VDD VSS BUF_X1 
XU557 n1432 n647 VDD VSS BUF_X1 
XU558 n1437 n648 VDD VSS BUF_X1 
XU559 n1448 n649 VDD VSS BUF_X1 
XU560 n1459 n650 VDD VSS BUF_X1 
XU561 n1469 n651 VDD VSS BUF_X1 
XU562 n1468 n652 VDD VSS CLKBUF_X1 
XU563 n1475 n653 VDD VSS BUF_X1 
XU564 n1480 n654 VDD VSS BUF_X1 
XU565 n1488 n655 VDD VSS INV_X1 
XU566 n655 n656 VDD VSS INV_X32 
XU567 n1496 n657 VDD VSS BUF_X1 
XU568 n1501 n658 VDD VSS BUF_X1 
XU569 n1506 n659 VDD VSS BUF_X1 
XU570 n1511 n660 VDD VSS INV_X1 
XU571 n660 n661 VDD VSS INV_X8 
XU572 n1516 n662 VDD VSS BUF_X1 
XU573 n1521 n663 VDD VSS BUF_X1 
XU574 n1526 n664 VDD VSS INV_X1 
XU575 n664 n665 VDD VSS INV_X16 
XU576 n1531 n666 VDD VSS BUF_X1 
XU577 n181 n667 VDD VSS CLKBUF_X1 
XU578 n1542 n668 VDD VSS BUF_X1 
XU579 n1547 n669 VDD VSS BUF_X1 
XU580 n1552 n670 VDD VSS INV_X1 
XU581 n670 n671 VDD VSS INV_X8 
XU582 n1575 n672 VDD VSS BUF_X1 
XU583 n1574 n673 VDD VSS CLKBUF_X1 
XU584 n1592 n674 VDD VSS BUF_X1 
XU585 n1597 n675 VDD VSS BUF_X1 
XU586 n1602 n676 VDD VSS INV_X1 
XU587 n676 n677 VDD VSS INV_X8 
XU588 n1611 n678 VDD VSS BUF_X1 
XU589 n1618 n679 VDD VSS BUF_X1 
XU590 n1623 n680 VDD VSS BUF_X1 
XU591 n1639 n681 VDD VSS BUF_X1 
XU592 n1638 n682 VDD VSS CLKBUF_X1 
XU593 n1651 n683 VDD VSS BUF_X1 
XU594 n1656 n684 VDD VSS BUF_X1 
XU595 n1661 n685 VDD VSS BUF_X1 
XU596 n1666 n686 VDD VSS BUF_X1 
XU597 n1671 n687 VDD VSS BUF_X1 
XU598 n1675 n688 VDD VSS BUF_X1 
XU599 n1674 n689 VDD VSS CLKBUF_X1 
XU600 n1678 n690 VDD VSS BUF_X1 
XU601 n1677 n691 VDD VSS CLKBUF_X1 
XU602 n1686 n692 VDD VSS BUF_X1 
XU603 n1697 n693 VDD VSS BUF_X1 
XU604 n1702 n694 VDD VSS BUF_X1 
XU605 n1713 n695 VDD VSS BUF_X1 
XU606 n1716 n696 VDD VSS CLKBUF_X1 
XU607 n1728 n697 VDD VSS BUF_X1 
XU608 n54 n698 VDD VSS CLKBUF_X1 
XU609 n1727 n699 VDD VSS CLKBUF_X1 
XU610 n33 n700 VDD VSS BUF_X1 
XU611 n26 n701 VDD VSS BUF_X1 
XU612 n1755 n702 VDD VSS BUF_X1 
XU613 n19 n703 VDD VSS BUF_X1 
XU614 n1760 n704 VDD VSS CLKBUF_X1 
XU615 n1762 n705 VDD VSS BUF_X1 
XU616 n1761 n706 VDD VSS CLKBUF_X1 
XU617 n1770 n707 VDD VSS BUF_X1 
XU618 n1781 n708 VDD VSS BUF_X1 
XU619 n1786 n709 VDD VSS BUF_X1 
XU620 n1795 n710 VDD VSS BUF_X1 
XU621 n1802 n711 VDD VSS CLKBUF_X1 
XU622 n1813 n712 VDD VSS BUF_X1 
XU623 n1818 n713 VDD VSS BUF_X1 
XU624 n1823 n714 VDD VSS BUF_X1 
XU625 n1828 n715 VDD VSS BUF_X1 
XU626 n1833 n716 VDD VSS BUF_X1 
XU627 n1844 n717 VDD VSS CLKBUF_X1 
XU628 n1852 n718 VDD VSS BUF_X1 
XU629 n49 n719 VDD VSS CLKBUF_X1 
XU630 n1859 n720 VDD VSS BUF_X1 
XU631 n1868 n721 VDD VSS BUF_X1 
XU632 n1875 n722 VDD VSS BUF_X1 
XU633 n1878 n723 VDD VSS CLKBUF_X1 
XU634 n1885 n724 VDD VSS BUF_X1 
XU635 n1884 n725 VDD VSS CLKBUF_X1 
XU636 n45 n726 VDD VSS BUF_X1 
XU637 n38 n727 VDD VSS BUF_X1 
XU638 n1904 n728 VDD VSS BUF_X1 
XU639 n31 n729 VDD VSS BUF_X1 
XU640 n1911 n730 VDD VSS BUF_X1 
XU641 n1916 n731 VDD VSS BUF_X1 
XU642 n17 n732 VDD VSS BUF_X1 
XU643 n1921 n733 VDD VSS CLKBUF_X1 
XU644 n1930 n734 VDD VSS BUF_X1 
XU645 n123 n735 VDD VSS CLKBUF_X1 
XU646 n1929 n736 VDD VSS CLKBUF_X1 
XU647 n1942 n737 VDD VSS INV_X1 
XU648 n737 n738 VDD VSS INV_X4 
XU649 n1947 n739 VDD VSS BUF_X1 
XU650 n1958 n740 VDD VSS BUF_X1 
XU651 n1963 n741 VDD VSS BUF_X1 
XU652 n1968 n742 VDD VSS CLKBUF_X1 
XU653 n1972 n743 VDD VSS INV_X1 
XU654 n743 n744 VDD VSS INV_X32 
XU655 n1985 n745 VDD VSS BUF_X1 
XU656 n1990 n746 VDD VSS BUF_X1 
XU657 n1995 n747 VDD VSS BUF_X1 
XU658 n2012 n748 VDD VSS BUF_X1 
XU659 n752 n749 VDD VSS CLKBUF_X1 
XU660 n749 n750 VDD VSS INV_X32 
XU661 n750 n751 VDD VSS INV_X1 
XU662 n402 n752 VDD VSS INV_X1 
XU663 n751 n753 VDD VSS INV_X32 
XU664 n757 n754 VDD VSS CLKBUF_X1 
XU665 n754 n755 VDD VSS INV_X32 
XU666 n755 n756 VDD VSS INV_X1 
XU667 n389 n757 VDD VSS INV_X1 
XU668 n756 n758 VDD VSS INV_X32 
XU669 n762 n759 VDD VSS CLKBUF_X1 
XU670 n759 n760 VDD VSS INV_X32 
XU671 n760 n761 VDD VSS INV_X1 
XU672 n376 n762 VDD VSS INV_X1 
XU673 n761 n763 VDD VSS INV_X32 
XU674 n769 n764 VDD VSS INV_X1 
XU675 n764 n765 VDD VSS INV_X32 
XU676 n768 n766 VDD VSS INV_X32 
XU677 n766 n767 VDD VSS INV_X1 
XU678 n421 n768 VDD VSS INV_X1 
XU679 n767 n769 VDD VSS INV_X32 
XU680 n408 n770 VDD VSS INV_X1 
XU681 n770 n771 VDD VSS INV_X32 
XU682 n771 n772 VDD VSS INV_X1 
XU683 n562 n773 VDD VSS INV_X32 
XU684 n159 n774 VDD VSS CLKBUF_X1 
XU685 n778 n775 VDD VSS CLKBUF_X1 
XU686 n775 n776 VDD VSS INV_X32 
XU687 n776 n777 VDD VSS INV_X1 
XU688 n395 n778 VDD VSS INV_X1 
XU689 n777 n779 VDD VSS INV_X32 
XU690 n783 n780 VDD VSS CLKBUF_X1 
XU691 n382 n781 VDD VSS INV_X1 
XU692 n781 n782 VDD VSS INV_X32 
XU693 n782 n783 VDD VSS INV_X1 
XU694 n780 n784 VDD VSS INV_X32 
XU695 n788 n785 VDD VSS CLKBUF_X1 
XU696 n785 n786 VDD VSS INV_X32 
XU697 n566 n787 VDD VSS INV_X1 
XU698 n427 n788 VDD VSS INV_X1 
XU699 n787 n789 VDD VSS INV_X32 
XU700 n793 n790 VDD VSS CLKBUF_X1 
XU701 n790 n791 VDD VSS INV_X32 
XU702 n568 n792 VDD VSS INV_X1 
XU703 n414 n793 VDD VSS INV_X1 
XU704 n792 n794 VDD VSS INV_X32 
XU705 n798 n795 VDD VSS CLKBUF_X1 
XU706 n795 n796 VDD VSS INV_X32 
XU707 n796 n797 VDD VSS INV_X1 
XU708 n401 n798 VDD VSS INV_X1 
XU709 n797 n799 VDD VSS INV_X32 
XU710 n803 n800 VDD VSS CLKBUF_X1 
XU711 n388 n801 VDD VSS INV_X1 
XU712 n801 n802 VDD VSS INV_X32 
XU713 n802 n803 VDD VSS INV_X1 
XU714 n800 n804 VDD VSS INV_X32 
XU715 n8 n805 VDD VSS INV_X1 
XU716 n805 n806 VDD VSS INV_X32 
XU717 n233 n807 VDD VSS INV_X1 
XU718 n807 n808 VDD VSS INV_X32 
XU719 N3091 n809 VDD VSS INV_X1 
XU720 n809 n810 VDD VSS INV_X32 
XU721 n816 n811 VDD VSS INV_X1 
XU723 n235 n813 VDD VSS INV_X1 
XU724 n813 n814 VDD VSS INV_X32 
XU725 N3081 n815 VDD VSS INV_X1 
XU726 n815 n816 VDD VSS INV_X32 
XU727 n822 n817 VDD VSS INV_X1 
XU728 n817 n818 VDD VSS INV_X16 
XU729 n237 n819 VDD VSS INV_X1 
XU730 n819 n820 VDD VSS INV_X32 
XU731 N3071 n821 VDD VSS INV_X1 
XU732 n821 n822 VDD VSS INV_X32 
XU733 n828 n823 VDD VSS INV_X1 
XU734 n823 n824 VDD VSS INV_X8 
XU735 n239 n825 VDD VSS INV_X1 
XU736 n825 n826 VDD VSS INV_X32 
XU737 N3061 n827 VDD VSS INV_X1 
XU738 n827 n828 VDD VSS INV_X32 
XU739 n834 n829 VDD VSS INV_X1 
XU740 n829 n830 VDD VSS INV_X8 
XU741 n241 n831 VDD VSS INV_X1 
XU742 n831 n832 VDD VSS INV_X32 
XU743 N3051 n833 VDD VSS INV_X1 
XU744 n833 n834 VDD VSS INV_X32 
XU745 n840 n835 VDD VSS INV_X1 
XU746 n835 n836 VDD VSS INV_X32 
XU747 n243 n837 VDD VSS INV_X1 
XU748 n837 n838 VDD VSS INV_X32 
XU749 N3041 n839 VDD VSS INV_X1 
XU750 n839 n840 VDD VSS INV_X32 
XU751 n845 n841 VDD VSS CLKBUF_X1 
XU752 n245 n842 VDD VSS INV_X1 
XU753 n842 n843 VDD VSS INV_X32 
XU754 N303 n844 VDD VSS INV_X1 
XU755 n844 n845 VDD VSS INV_X32 
XU756 n850 n846 VDD VSS BUF_X1 
XU757 n2470 n847 VDD VSS INV_X1 
XU758 n847 n848 VDD VSS INV_X32 
XU759 N302 n849 VDD VSS INV_X1 
XU760 n849 n850 VDD VSS INV_X32 
XU761 n856 n851 VDD VSS INV_X1 
XU762 n851 n852 VDD VSS INV_X32 
XU763 n2490 n853 VDD VSS INV_X1 
XU764 n853 n854 VDD VSS INV_X32 
XU765 N301 n855 VDD VSS INV_X1 
XU766 n855 n856 VDD VSS INV_X32 
XU767 n862 n857 VDD VSS INV_X1 
XU768 n857 n858 VDD VSS INV_X32 
XU769 n2510 n859 VDD VSS INV_X1 
XU770 n859 n860 VDD VSS INV_X32 
XU771 N300 n861 VDD VSS INV_X1 
XU772 n861 n862 VDD VSS INV_X32 
XU773 n866 n863 VDD VSS INV_X1 
XU774 n863 n864 VDD VSS INV_X16 
XU775 N299 n865 VDD VSS INV_X1 
XU776 n865 n866 VDD VSS INV_X32 
XU777 n2530 n867 VDD VSS INV_X1 
XU778 n867 n868 VDD VSS INV_X32 
XU779 n872 n869 VDD VSS INV_X1 
XU780 n869 n870 VDD VSS INV_X16 
XU781 N298 n871 VDD VSS INV_X1 
XU782 n871 n872 VDD VSS INV_X32 
XU783 n25500 n873 VDD VSS INV_X1 
XU784 n873 n874 VDD VSS INV_X32 
XU785 n880 n875 VDD VSS INV_X1 
XU786 n875 n876 VDD VSS INV_X8 
XU787 n25700 n877 VDD VSS INV_X1 
XU788 n877 n878 VDD VSS INV_X32 
XU789 N297 n879 VDD VSS INV_X1 
XU790 n879 n880 VDD VSS INV_X32 
XU791 n884 n881 VDD VSS INV_X1 
XU792 n881 n882 VDD VSS INV_X16 
XU793 N296 n883 VDD VSS INV_X1 
XU794 n883 n884 VDD VSS INV_X32 
XU795 n25900 n885 VDD VSS INV_X1 
XU796 n885 n886 VDD VSS INV_X32 
XU797 n892 n887 VDD VSS INV_X1 
XU798 n887 n888 VDD VSS INV_X8 
XU799 n26100 n889 VDD VSS INV_X1 
XU800 n889 n890 VDD VSS INV_X32 
XU801 N295 n891 VDD VSS INV_X1 
XU802 n891 n892 VDD VSS INV_X32 
XU803 n898 n893 VDD VSS INV_X1 
XU804 n893 n894 VDD VSS INV_X16 
XU805 n2630 n895 VDD VSS INV_X1 
XU806 n895 n896 VDD VSS INV_X32 
XU807 N294 n897 VDD VSS INV_X1 
XU808 n897 n898 VDD VSS INV_X32 
XU809 n904 n899 VDD VSS INV_X1 
XU810 n899 n900 VDD VSS INV_X8 
XU811 n2650 n901 VDD VSS INV_X1 
XU812 n901 n902 VDD VSS INV_X32 
XU813 N293 n903 VDD VSS INV_X1 
XU814 n903 n904 VDD VSS INV_X32 
XU815 n910 n905 VDD VSS INV_X1 
XU816 n905 n906 VDD VSS INV_X16 
XU817 n2670 n907 VDD VSS INV_X1 
XU818 n907 n908 VDD VSS INV_X32 
XU819 N292 n909 VDD VSS INV_X1 
XU820 n909 n910 VDD VSS INV_X32 
XU821 n916 n911 VDD VSS INV_X1 
XU822 n2690 n913 VDD VSS INV_X1 
XU823 n913 n914 VDD VSS INV_X32 
XU824 N291 n915 VDD VSS INV_X1 
XU825 n915 n916 VDD VSS INV_X32 
XU826 n922 n917 VDD VSS INV_X1 
XU827 n917 n918 VDD VSS INV_X8 
XU828 n2710 n919 VDD VSS INV_X1 
XU829 n919 n920 VDD VSS INV_X32 
XU830 N290 n921 VDD VSS INV_X1 
XU831 n921 n922 VDD VSS INV_X32 
XU832 n928 n923 VDD VSS INV_X1 
XU833 n923 n924 VDD VSS INV_X16 
XU834 n2730 n925 VDD VSS INV_X1 
XU835 n925 n926 VDD VSS INV_X32 
XU836 N289 n927 VDD VSS INV_X1 
XU837 n927 n928 VDD VSS INV_X32 
XU838 n934 n929 VDD VSS INV_X1 
XU839 n929 n930 VDD VSS INV_X32 
XU840 n2750 n931 VDD VSS INV_X1 
XU841 n931 n932 VDD VSS INV_X32 
XU842 N288 n933 VDD VSS INV_X1 
XU843 n933 n934 VDD VSS INV_X32 
XU844 N287 n935 VDD VSS INV_X1 
XU845 n935 n936 VDD VSS INV_X32 
XU846 n2770 n937 VDD VSS INV_X1 
XU847 n937 n938 VDD VSS INV_X32 
XU848 n2790 n939 VDD VSS INV_X1 
XU849 n939 n940 VDD VSS INV_X32 
XU850 N286 n941 VDD VSS INV_X1 
XU851 n941 n942 VDD VSS INV_X32 
XU852 n948 n943 VDD VSS INV_X1 
XU853 n943 n944 VDD VSS INV_X16 
XU854 n2810 n945 VDD VSS INV_X1 
XU855 n945 n946 VDD VSS INV_X32 
XU856 N285 n947 VDD VSS INV_X1 
XU857 n947 n948 VDD VSS INV_X32 
XU858 n954 n949 VDD VSS INV_X1 
XU859 n949 n950 VDD VSS INV_X16 
XU860 n2830 n951 VDD VSS INV_X1 
XU861 n951 n952 VDD VSS INV_X32 
XU862 N284 n953 VDD VSS INV_X1 
XU863 n953 n954 VDD VSS INV_X32 
XU864 n960 n955 VDD VSS INV_X1 
XU865 n955 n956 VDD VSS INV_X8 
XU866 n2850 n957 VDD VSS INV_X1 
XU867 n957 n958 VDD VSS INV_X32 
XU868 N283 n959 VDD VSS INV_X1 
XU869 n959 n960 VDD VSS INV_X32 
XU870 n966 n961 VDD VSS INV_X1 
XU871 n2870 n963 VDD VSS INV_X1 
XU872 n963 n964 VDD VSS INV_X32 
XU873 N282 n965 VDD VSS INV_X1 
XU874 n965 n966 VDD VSS INV_X32 
XU875 n972 n967 VDD VSS INV_X1 
XU876 n967 n968 VDD VSS INV_X32 
XU877 n2890 n969 VDD VSS INV_X1 
XU878 n969 n970 VDD VSS INV_X32 
XU879 N281 n971 VDD VSS INV_X1 
XU880 n971 n972 VDD VSS INV_X32 
XU881 n975 n973 VDD VSS BUF_X1 
XU882 N280 n974 VDD VSS INV_X1 
XU883 n974 n975 VDD VSS INV_X32 
XU884 n2910 n976 VDD VSS INV_X1 
XU885 n976 n977 VDD VSS INV_X32 
XU886 n983 n978 VDD VSS INV_X1 
XU887 n978 n979 VDD VSS INV_X16 
XU888 n2930 n980 VDD VSS INV_X1 
XU889 n980 n981 VDD VSS INV_X32 
XU890 N279 n982 VDD VSS INV_X1 
XU891 n982 n983 VDD VSS INV_X32 
XU892 n989 n984 VDD VSS INV_X1 
XU893 n984 n985 VDD VSS INV_X16 
XU894 n2950 n986 VDD VSS INV_X1 
XU895 n986 n987 VDD VSS INV_X32 
XU896 N278 n988 VDD VSS INV_X1 
XU897 n988 n989 VDD VSS INV_X32 
XU898 n995 n990 VDD VSS INV_X1 
XU899 n2970 n992 VDD VSS INV_X1 
XU900 n992 n993 VDD VSS INV_X32 
XU901 N277 n994 VDD VSS INV_X1 
XU902 n994 n995 VDD VSS INV_X32 
XU903 n1001 n996 VDD VSS INV_X1 
XU904 n996 n997 VDD VSS INV_X16 
XU905 n2990 n998 VDD VSS INV_X1 
XU906 n998 n999 VDD VSS INV_X32 
XU907 N276 n1000 VDD VSS INV_X1 
XU908 n1000 n1001 VDD VSS INV_X32 
XU909 n1005 n1002 VDD VSS INV_X1 
XU910 n1002 n1003 VDD VSS INV_X16 
XU911 N275 n1004 VDD VSS INV_X1 
XU912 n1004 n1005 VDD VSS INV_X32 
XU913 n3010 n1006 VDD VSS INV_X1 
XU914 n1006 n1007 VDD VSS INV_X32 
XU915 N274 n1008 VDD VSS INV_X1 
XU916 n1008 n1009 VDD VSS INV_X32 
XU917 n3030 n1010 VDD VSS INV_X1 
XU918 n1010 n1011 VDD VSS INV_X32 
XU919 N273 n1013 VDD VSS INV_X1 
XU920 n1013 n1014 VDD VSS INV_X32 
XU921 n1012 n1015 VDD VSS INV_X1 
XU922 n1015 n1016 VDD VSS INV_X32 
XU923 n1022 n1017 VDD VSS INV_X1 
XU924 n1017 n1018 VDD VSS INV_X16 
XU925 n3070 n1019 VDD VSS INV_X1 
XU926 n1019 n1020 VDD VSS INV_X32 
XU927 N272 n1021 VDD VSS INV_X1 
XU928 n1021 n1022 VDD VSS INV_X32 
XU929 n1027 n1023 VDD VSS BUF_X1 
XU930 n3090 n1024 VDD VSS INV_X1 
XU931 n1024 n1025 VDD VSS INV_X32 
XU932 N271 n1026 VDD VSS INV_X1 
XU933 n1026 n1027 VDD VSS INV_X32 
XU934 n1033 n1028 VDD VSS INV_X1 
XU935 n1028 n1029 VDD VSS INV_X16 
XU936 n311 n1030 VDD VSS INV_X1 
XU937 n1030 n1031 VDD VSS INV_X32 
XU938 N270 n1032 VDD VSS INV_X1 
XU939 n1032 n1033 VDD VSS INV_X32 
XU940 n1039 n1034 VDD VSS INV_X1 
XU941 n1034 n1035 VDD VSS INV_X32 
XU942 n313 n1036 VDD VSS INV_X1 
XU943 n1036 n1037 VDD VSS INV_X32 
XU944 N269 n1038 VDD VSS INV_X1 
XU945 n1038 n1039 VDD VSS INV_X32 
XU946 n1041 n1040 VDD VSS CLKBUF_X1 
XU947 n315 n1041 VDD VSS INV_X1 
XU948 n1040 n1042 VDD VSS INV_X32 
XU949 N268 n1043 VDD VSS INV_X1 
XU950 n1043 n1044 VDD VSS INV_X32 
XU951 n1049 n1045 VDD VSS BUF_X1 
XU952 n317 n1046 VDD VSS INV_X1 
XU953 n1046 n1047 VDD VSS INV_X32 
XU954 N267 n1048 VDD VSS INV_X1 
XU955 n1048 n1049 VDD VSS INV_X32 
XU956 n1055 n1050 VDD VSS INV_X1 
XU957 n1050 n1051 VDD VSS INV_X16 
XU958 n319 n1052 VDD VSS INV_X1 
XU959 n1052 n1053 VDD VSS INV_X32 
XU960 N266 n1054 VDD VSS INV_X1 
XU961 n1054 n1055 VDD VSS INV_X32 
XU962 n1060 n1056 VDD VSS BUF_X1 
XU963 n321 n1057 VDD VSS INV_X1 
XU964 n1057 n1058 VDD VSS INV_X32 
XU965 N265 n1059 VDD VSS INV_X1 
XU966 n1059 n1060 VDD VSS INV_X32 
XU967 n1062 n1061 VDD VSS CLKBUF_X1 
XU968 n323 n1062 VDD VSS INV_X1 
XU969 n1061 n1063 VDD VSS INV_X32 
XU970 N264 n1064 VDD VSS INV_X1 
XU971 n1064 n1065 VDD VSS INV_X32 
XU972 n1070 n1066 VDD VSS BUF_X1 
XU973 n325 n1067 VDD VSS INV_X1 
XU974 n1067 n1068 VDD VSS INV_X32 
XU975 N263 n1069 VDD VSS INV_X1 
XU976 n1069 n1070 VDD VSS INV_X32 
XU977 n1075 n1071 VDD VSS BUF_X1 
XU978 n327 n1072 VDD VSS INV_X1 
XU979 n1072 n1073 VDD VSS INV_X32 
XU980 N262 n1074 VDD VSS INV_X1 
XU981 n1074 n1075 VDD VSS INV_X32 
XU982 n1078 n1076 VDD VSS BUF_X1 
XU983 N2610 n1077 VDD VSS INV_X1 
XU984 n1077 n1078 VDD VSS INV_X32 
XU985 n329 n1079 VDD VSS INV_X1 
XU986 n1079 n1080 VDD VSS INV_X32 
XU987 n1084 n1081 VDD VSS INV_X1 
XU988 n1081 n1082 VDD VSS INV_X32 
XU989 N2600 n1083 VDD VSS INV_X1 
XU990 n1083 n1084 VDD VSS INV_X32 
XU991 n1088 n1085 VDD VSS INV_X1 
XU992 n1085 n1086 VDD VSS INV_X32 
XU993 N2590 n1087 VDD VSS INV_X1 
XU994 n1087 n1088 VDD VSS INV_X32 
XU995 n335 n1089 VDD VSS INV_X1 
XU996 n1089 n1090 VDD VSS INV_X32 
XU997 N2580 n1091 VDD VSS INV_X1 
XU998 n1091 n1092 VDD VSS INV_X32 
XU999 n1097 n1093 VDD VSS BUF_X1 
XU1000 n337 n1094 VDD VSS INV_X1 
XU1001 n1094 n1095 VDD VSS INV_X32 
XU1002 N2570 n1096 VDD VSS INV_X1 
XU1003 n1096 n1097 VDD VSS INV_X32 
XU1004 n1102 n1098 VDD VSS BUF_X1 
XU1005 n339 n1099 VDD VSS INV_X1 
XU1006 n1099 n1100 VDD VSS INV_X32 
XU1007 N2560 n1101 VDD VSS INV_X1 
XU1008 n1101 n1102 VDD VSS INV_X32 
XU1009 n1104 n1103 VDD VSS CLKBUF_X1 
XU1010 n341 n1104 VDD VSS INV_X1 
XU1011 n1103 n1105 VDD VSS INV_X32 
XU1012 N2550 n1106 VDD VSS INV_X1 
XU1013 n1106 n1107 VDD VSS INV_X32 
XU1014 n1108 n1109 VDD VSS INV_X1 
XU1015 n1109 n1110 VDD VSS INV_X32 
XU1016 N2540 n1111 VDD VSS INV_X1 
XU1017 n1111 n1112 VDD VSS INV_X32 
XU1018 n1114 n1113 VDD VSS CLKBUF_X1 
XU1019 n346 n1114 VDD VSS INV_X1 
XU1020 n1113 n1115 VDD VSS INV_X32 
XU1021 N253 n1116 VDD VSS INV_X1 
XU1022 n1116 n1117 VDD VSS INV_X32 
XU1023 n1122 n1118 VDD VSS BUF_X1 
XU1024 n349 n1119 VDD VSS INV_X1 
XU1025 n1119 n1120 VDD VSS INV_X32 
XU1026 N2520 n1121 VDD VSS INV_X1 
XU1027 n1121 n1122 VDD VSS INV_X32 
XU1028 n352 n1123 VDD VSS INV_X1 
XU1029 n1123 n1124 VDD VSS INV_X32 
XU1030 N251 n1125 VDD VSS INV_X1 
XU1031 n1125 n1126 VDD VSS INV_X32 
XU1032 n1131 n1127 VDD VSS BUF_X1 
XU1033 n356 n1128 VDD VSS INV_X1 
XU1034 n1128 n1129 VDD VSS INV_X32 
XU1035 N2500 n1130 VDD VSS INV_X1 
XU1036 n1130 n1131 VDD VSS INV_X32 
XU1037 n1136 n1132 VDD VSS BUF_X1 
XU1038 n360 n1133 VDD VSS INV_X1 
XU1039 n1133 n1134 VDD VSS INV_X32 
XU1040 N249 n1135 VDD VSS INV_X1 
XU1041 n1135 n1136 VDD VSS INV_X32 
XU1042 n1141 n1137 VDD VSS BUF_X1 
XU1043 n364 n1138 VDD VSS INV_X1 
XU1044 n1138 n1139 VDD VSS INV_X32 
XU1045 N2480 n1140 VDD VSS INV_X1 
XU1046 n1140 n1141 VDD VSS INV_X32 
XU1047 n1146 n1142 VDD VSS BUF_X1 
XU1048 n368 n1143 VDD VSS INV_X1 
XU1049 n1143 n1144 VDD VSS INV_X32 
XU1050 N247 n1145 VDD VSS INV_X1 
XU1051 n1145 n1146 VDD VSS INV_X32 
XU1052 n372 n1147 VDD VSS INV_X1 
XU1053 n1147 n1148 VDD VSS INV_X32 
XU1054 N2460 n1149 VDD VSS INV_X1 
XU1055 n1149 n1150 VDD VSS INV_X32 
XU1056 n164 n1151 VDD VSS INV_X32 
XU1057 n1151 n1152 VDD VSS INV_X1 
XU1058 n1156 n1153 VDD VSS CLKBUF_X1 
XU1059 n1153 n1154 VDD VSS INV_X32 
XU1060 n1154 n1155 VDD VSS INV_X1 
XU1061 n470 n1156 VDD VSS INV_X1 
XU1062 n1155 n1157 VDD VSS INV_X32 
XU1063 n1161 n1158 VDD VSS CLKBUF_X1 
XU1064 n1158 n1159 VDD VSS INV_X32 
XU1065 n579 n1160 VDD VSS INV_X1 
XU1066 n446 n1161 VDD VSS INV_X1 
XU1067 n1160 n1162 VDD VSS INV_X32 
XU1068 n1164 n1163 VDD VSS CLKBUF_X1 
XU1069 n480 n1164 VDD VSS INV_X1 
XU1070 n1163 n1165 VDD VSS INV_X32 
XU1071 n1165 n1166 VDD VSS INV_X1 
XU1072 n1166 n1167 VDD VSS INV_X32 
XU1073 n1173 n1168 VDD VSS INV_X1 
XU1074 n1168 n1169 VDD VSS INV_X32 
XU1075 n1172 n1170 VDD VSS INV_X32 
XU1076 n1170 n1171 VDD VSS INV_X1 
XU1077 n456 n1172 VDD VSS INV_X1 
XU1078 n1171 n1173 VDD VSS INV_X32 
XU1079 n1177 n1174 VDD VSS CLKBUF_X1 
XU1080 n1174 n1175 VDD VSS INV_X32 
XU1081 n1175 n1176 VDD VSS INV_X1 
XU1082 n495 n1177 VDD VSS INV_X1 
XU1083 n1176 n1178 VDD VSS INV_X32 
XU1084 n1182 n1179 VDD VSS CLKBUF_X1 
XU1085 n1179 n1180 VDD VSS INV_X32 
XU1086 n1180 n1181 VDD VSS INV_X1 
XU1087 n471 n1182 VDD VSS INV_X1 
XU1088 n1181 n1183 VDD VSS INV_X32 
XU1089 n1187 n1184 VDD VSS CLKBUF_X1 
XU1090 n447 n1185 VDD VSS INV_X1 
XU1091 n1185 n1186 VDD VSS INV_X32 
XU1092 n585 n1187 VDD VSS INV_X1 
XU1093 n1184 n1188 VDD VSS INV_X32 
XU1094 n1190 n1189 VDD VSS CLKBUF_X1 
XU1095 n481 n1190 VDD VSS INV_X1 
XU1096 n1189 n1191 VDD VSS INV_X32 
XU1097 n1191 n1192 VDD VSS INV_X1 
XU1098 n1192 n1193 VDD VSS INV_X32 
XU1099 n1197 n1194 VDD VSS CLKBUF_X1 
XU1100 n457 n1195 VDD VSS INV_X1 
XU1101 n1195 n1196 VDD VSS INV_X32 
XU1102 n1196 n1197 VDD VSS INV_X1 
XU1103 n1194 n1198 VDD VSS INV_X32 
XU1104 n1202 n1199 VDD VSS CLKBUF_X1 
XU1105 n1199 n1200 VDD VSS INV_X32 
XU1106 n1200 n1201 VDD VSS INV_X1 
XU1107 n491 n1202 VDD VSS INV_X1 
XU1108 n1201 n1203 VDD VSS INV_X32 
XU1109 n1207 n1204 VDD VSS CLKBUF_X1 
XU1110 n1204 n1205 VDD VSS INV_X32 
XU1111 n1205 n1206 VDD VSS INV_X1 
XU1112 n467 n1207 VDD VSS INV_X1 
XU1113 n1206 n1208 VDD VSS INV_X32 
XU1114 n1212 n1209 VDD VSS CLKBUF_X1 
XU1115 n1209 n1210 VDD VSS INV_X32 
XU1116 n1210 n1211 VDD VSS INV_X1 
XU1117 n443 n1212 VDD VSS INV_X1 
XU1118 n1211 n1213 VDD VSS INV_X32 
XU1119 n1217 n1214 VDD VSS CLKBUF_X1 
XU1120 n1214 n1215 VDD VSS INV_X32 
XU1121 n1215 n1216 VDD VSS INV_X1 
XU1122 n477 n1217 VDD VSS INV_X1 
XU1123 n1216 n1218 VDD VSS INV_X32 
XU1124 n1222 n1219 VDD VSS CLKBUF_X1 
XU1125 n1219 n1220 VDD VSS INV_X32 
XU1126 n595 n1221 VDD VSS INV_X1 
XU1127 n453 n1222 VDD VSS INV_X1 
XU1128 n1221 n1223 VDD VSS INV_X32 
XU1129 n1225 n1224 VDD VSS CLKBUF_X1 
XU1130 n487 n1225 VDD VSS INV_X1 
XU1131 n1224 n1226 VDD VSS INV_X32 
XU1132 n1226 n1227 VDD VSS INV_X1 
XU1133 n1227 n1228 VDD VSS INV_X32 
XU1134 n1230 n1229 VDD VSS CLKBUF_X1 
XU1135 n463 n1230 VDD VSS INV_X1 
XU1136 n1229 n1231 VDD VSS INV_X32 
XU1137 n1231 n1232 VDD VSS INV_X1 
XU1138 n1232 n1233 VDD VSS INV_X32 
XU1139 n1238 n1234 VDD VSS BUF_X1 
XU1140 n1237 n1235 VDD VSS INV_X32 
XU1141 n1235 n1236 VDD VSS INV_X1 
XU1142 n439 n1237 VDD VSS INV_X1 
XU1143 n1236 n1238 VDD VSS INV_X32 
XU1144 n1242 n1239 VDD VSS CLKBUF_X1 
XU1145 n1239 n1240 VDD VSS INV_X32 
XU1146 n1240 n1241 VDD VSS INV_X1 
XU1147 n473 n1242 VDD VSS INV_X1 
XU1148 n1241 n1243 VDD VSS INV_X32 
XU1149 n1247 n1244 VDD VSS CLKBUF_X1 
XU1150 n449 n1245 VDD VSS INV_X1 
XU1151 n1245 n1246 VDD VSS INV_X32 
XU1152 n600 n1247 VDD VSS INV_X1 
XU1153 n1244 n1248 VDD VSS INV_X32 
XU1154 n1254 n1249 VDD VSS INV_X1 
XU1155 n1249 n1250 VDD VSS INV_X32 
XU1156 n488 n1251 VDD VSS INV_X1 
XU1157 n1251 n1252 VDD VSS INV_X32 
XU1158 n1252 n1253 VDD VSS INV_X1 
XU1159 n1253 n1254 VDD VSS INV_X32 
XU1160 n1258 n1255 VDD VSS CLKBUF_X1 
XU1161 n1255 n1256 VDD VSS INV_X32 
XU1162 n1256 n1257 VDD VSS INV_X1 
XU1163 n464 n1258 VDD VSS INV_X1 
XU1164 n1257 n1259 VDD VSS INV_X32 
XU1165 n1265 n1260 VDD VSS INV_X1 
XU1166 n1260 n1261 VDD VSS INV_X32 
XU1167 n440 n1262 VDD VSS INV_X1 
XU1168 n1262 n1263 VDD VSS INV_X32 
XU1169 n1263 n1264 VDD VSS INV_X1 
XU1170 n1264 n1265 VDD VSS INV_X32 
XU1171 n1269 n1266 VDD VSS CLKBUF_X1 
XU1172 n483 n1267 VDD VSS INV_X1 
XU1173 n1267 n1268 VDD VSS INV_X32 
XU1174 n603 n1269 VDD VSS INV_X1 
XU1175 n1266 n1270 VDD VSS INV_X32 
XU1176 n1272 n1271 VDD VSS CLKBUF_X1 
XU1177 n459 n1272 VDD VSS INV_X1 
XU1178 n1271 n1273 VDD VSS INV_X32 
XU1179 n1273 n1274 VDD VSS INV_X1 
XU1180 n1274 n1275 VDD VSS INV_X32 
XU1181 n1279 n1276 VDD VSS CLKBUF_X1 
XU1182 n1276 n1277 VDD VSS INV_X32 
XU1183 n1277 n1278 VDD VSS INV_X1 
XU1184 n435 n1279 VDD VSS INV_X1 
XU1185 n1278 n1280 VDD VSS INV_X32 
XU1186 n1282 n1281 VDD VSS CLKBUF_X1 
XU1187 n474 n1282 VDD VSS INV_X1 
XU1188 n1281 n1283 VDD VSS INV_X32 
XU1189 n1283 n1284 VDD VSS INV_X1 
XU1190 n1284 n1285 VDD VSS INV_X32 
XU1191 n1289 n1286 VDD VSS CLKBUF_X1 
XU1192 n450 n1287 VDD VSS INV_X1 
XU1193 n1287 n1288 VDD VSS INV_X32 
XU1194 n1288 n1289 VDD VSS INV_X1 
XU1195 n1286 n1290 VDD VSS INV_X32 
XU1196 n1294 n1291 VDD VSS CLKBUF_X1 
XU1197 n1291 n1292 VDD VSS INV_X32 
XU1198 n1292 n1293 VDD VSS INV_X1 
XU1199 n489 n1294 VDD VSS INV_X1 
XU1200 n1293 n1295 VDD VSS INV_X32 
XU1201 n610 n1296 VDD VSS INV_X32 
XU1202 n1296 n1297 VDD VSS INV_X1 
XU1203 n465 n1298 VDD VSS INV_X1 
XU1204 n1297 n1299 VDD VSS INV_X32 
XU1205 n92 n1300 VDD VSS BUF_X1 
XU1206 n1304 n1301 VDD VSS CLKBUF_X1 
XU1207 n441 n1302 VDD VSS INV_X1 
XU1208 n1302 n1303 VDD VSS INV_X32 
XU1209 n1303 n1304 VDD VSS INV_X1 
XU1210 n1301 n1305 VDD VSS INV_X32 
XU1211 n1308 n1306 VDD VSS CLKBUF_X1 
XU1212 n1309 n1307 VDD VSS INV_X32 
XU1213 n1307 n1308 VDD VSS INV_X1 
XU1214 n484 n1309 VDD VSS INV_X1 
XU1215 n1306 n1310 VDD VSS INV_X32 
XU1216 n1314 n1311 VDD VSS CLKBUF_X1 
XU1217 n1311 n1312 VDD VSS INV_X32 
XU1218 n1312 n1313 VDD VSS INV_X1 
XU1219 n460 n1314 VDD VSS INV_X1 
XU1220 n1313 n1315 VDD VSS INV_X32 
XU1221 n1319 n1316 VDD VSS CLKBUF_X1 
XU1222 n1316 n1317 VDD VSS INV_X32 
XU1223 n1317 n1318 VDD VSS INV_X1 
XU1224 n436 n1319 VDD VSS INV_X1 
XU1225 n1318 n1320 VDD VSS INV_X32 
XU1226 n1324 n1321 VDD VSS CLKBUF_X1 
XU1227 n475 n1322 VDD VSS INV_X1 
XU1228 n1322 n1323 VDD VSS INV_X32 
XU1229 n1323 n1324 VDD VSS INV_X1 
XU1230 n1321 n1325 VDD VSS INV_X32 
XU1231 n1329 n1326 VDD VSS CLKBUF_X1 
XU1232 n451 n1327 VDD VSS INV_X1 
XU1233 n1327 n1328 VDD VSS INV_X32 
XU1234 n618 n1329 VDD VSS INV_X1 
XU1235 n1326 n1330 VDD VSS INV_X32 
XU1236 n1334 n1331 VDD VSS CLKBUF_X1 
XU1237 n1331 n1332 VDD VSS INV_X32 
XU1238 n1332 n1333 VDD VSS INV_X1 
XU1239 n490 n1334 VDD VSS INV_X1 
XU1240 n1333 n1335 VDD VSS INV_X32 
XU1241 n1339 n1336 VDD VSS CLKBUF_X1 
XU1242 n1336 n1337 VDD VSS INV_X32 
XU1243 n1337 n1338 VDD VSS INV_X1 
XU1244 n466 n1339 VDD VSS INV_X1 
XU1245 n1338 n1340 VDD VSS INV_X32 
XU1246 n1344 n1341 VDD VSS CLKBUF_X1 
XU1247 n1341 n1342 VDD VSS INV_X32 
XU1248 n1342 n1343 VDD VSS INV_X1 
XU1249 n442 n1344 VDD VSS INV_X1 
XU1250 n1343 n1345 VDD VSS INV_X32 
XU1251 n1349 n1346 VDD VSS CLKBUF_X1 
XU1252 n1346 n1347 VDD VSS INV_X32 
XU1253 n631 n1348 VDD VSS INV_X1 
XU1254 n485 n1349 VDD VSS INV_X1 
XU1255 n1348 n1350 VDD VSS INV_X32 
XU1256 n1354 n1351 VDD VSS CLKBUF_X1 
XU1257 n461 n1352 VDD VSS INV_X1 
XU1258 n1352 n1353 VDD VSS INV_X32 
XU1259 n1353 n1354 VDD VSS INV_X1 
XU1260 n1351 n1355 VDD VSS INV_X32 
XU1261 n1359 n1356 VDD VSS CLKBUF_X1 
XU1262 n437 n1357 VDD VSS INV_X1 
XU1263 n1357 n1358 VDD VSS INV_X32 
XU1264 n1358 n1359 VDD VSS INV_X1 
XU1265 n1356 n1360 VDD VSS INV_X32 
XU1266 n1364 n1361 VDD VSS CLKBUF_X1 
XU1267 n476 n1362 VDD VSS INV_X1 
XU1268 n1362 n1363 VDD VSS INV_X32 
XU1269 n1363 n1364 VDD VSS INV_X1 
XU1270 n1361 n1365 VDD VSS INV_X32 
XU1271 n1367 n1366 VDD VSS CLKBUF_X1 
XU1272 n452 n1367 VDD VSS INV_X1 
XU1273 n1366 n1368 VDD VSS INV_X32 
XU1274 n1368 n1369 VDD VSS INV_X1 
XU1275 n1369 n1370 VDD VSS INV_X32 
XU1276 n1372 n1371 VDD VSS CLKBUF_X1 
XU1277 n637 n1372 VDD VSS INV_X1 
XU1278 n1371 n1373 VDD VSS INV_X32 
XU1279 n486 n1374 VDD VSS INV_X1 
XU1280 n1374 n1375 VDD VSS INV_X32 
XU1281 n1379 n1376 VDD VSS CLKBUF_X1 
XU1282 n462 n1377 VDD VSS INV_X1 
XU1283 n1377 n1378 VDD VSS INV_X32 
XU1284 n1378 n1379 VDD VSS INV_X1 
XU1285 n1376 n1380 VDD VSS INV_X32 
XU1286 n1383 n1381 VDD VSS CLKBUF_X1 
XU1287 n1384 n1382 VDD VSS INV_X32 
XU1288 n1382 n1383 VDD VSS INV_X1 
XU1289 n438 n1384 VDD VSS INV_X1 
XU1290 n1381 n1385 VDD VSS INV_X32 
XU1291 n1391 n1386 VDD VSS INV_X1 
XU1292 n1386 n1387 VDD VSS INV_X32 
XU1293 n1390 n1388 VDD VSS INV_X32 
XU1294 n1388 n1389 VDD VSS INV_X1 
XU1295 n433 n1390 VDD VSS INV_X1 
XU1296 n1389 n1391 VDD VSS INV_X32 
XU1297 n420 n1392 VDD VSS INV_X1 
XU1298 n1392 n1393 VDD VSS INV_X32 
XU1299 n1393 n1394 VDD VSS INV_X1 
XU1300 n1394 n1395 VDD VSS INV_X32 
XU1301 n171 n1396 VDD VSS CLKBUF_X1 
XU1302 n1398 n1397 VDD VSS CLKBUF_X1 
XU1303 n407 n1398 VDD VSS INV_X1 
XU1304 n1397 n1399 VDD VSS INV_X32 
XU1305 n1399 n1400 VDD VSS INV_X1 
XU1306 n1400 n1401 VDD VSS INV_X32 
XU1307 n644 n1402 VDD VSS INV_X32 
XU1308 n1402 n1403 VDD VSS INV_X1 
XU1309 n394 n1404 VDD VSS INV_X1 
XU1310 n1403 n1405 VDD VSS INV_X32 
XU1311 n145 n1406 VDD VSS BUF_X1 
XU1312 n1410 n1407 VDD VSS CLKBUF_X1 
XU1313 n1407 n1408 VDD VSS INV_X32 
XU1314 n1408 n1409 VDD VSS INV_X1 
XU1315 n381 n1410 VDD VSS INV_X1 
XU1316 n1409 n1411 VDD VSS INV_X32 
XU1317 n1416 n1412 VDD VSS BUF_X1 
XU1318 n1415 n1413 VDD VSS INV_X32 
XU1319 n1413 n1414 VDD VSS INV_X1 
XU1320 n426 n1415 VDD VSS INV_X1 
XU1321 n1414 n1416 VDD VSS INV_X32 
XU1322 n177 n1417 VDD VSS INV_X1 
XU1323 n1417 n1418 VDD VSS INV_X32 
XU1324 n413 n1419 VDD VSS INV_X1 
XU1325 n1419 n1420 VDD VSS INV_X32 
XU1326 n1420 n1421 VDD VSS INV_X1 
XU1327 n1421 n1422 VDD VSS INV_X32 
XU1328 n1424 n1423 VDD VSS CLKBUF_X1 
XU1329 n400 n1424 VDD VSS INV_X1 
XU1330 n1423 n1425 VDD VSS INV_X32 
XU1331 n1425 n1426 VDD VSS INV_X1 
XU1332 n1426 n1427 VDD VSS INV_X32 
XU1333 n1429 n1428 VDD VSS CLKBUF_X1 
XU1334 n387 n1429 VDD VSS INV_X1 
XU1335 n1428 n1430 VDD VSS INV_X32 
XU1336 n1430 n1431 VDD VSS INV_X1 
XU1337 n1431 n1432 VDD VSS INV_X32 
XU1338 n1436 n1433 VDD VSS CLKBUF_X1 
XU1339 n1433 n1434 VDD VSS INV_X32 
XU1340 n1434 n1435 VDD VSS INV_X1 
XU1341 n432 n1436 VDD VSS INV_X1 
XU1342 n1435 n1437 VDD VSS INV_X32 
XU1343 n1443 n1438 VDD VSS INV_X1 
XU1344 n1438 n1439 VDD VSS INV_X32 
XU1345 n1442 n1440 VDD VSS INV_X32 
XU1346 n1440 n1441 VDD VSS INV_X1 
XU1347 n419 n1442 VDD VSS INV_X1 
XU1348 n1441 n1443 VDD VSS INV_X32 
XU1349 n1447 n1444 VDD VSS CLKBUF_X1 
XU1350 n1444 n1445 VDD VSS INV_X32 
XU1351 n1445 n1446 VDD VSS INV_X1 
XU1352 n406 n1447 VDD VSS INV_X1 
XU1353 n1446 n1448 VDD VSS INV_X32 
XU1354 n1454 n1449 VDD VSS INV_X1 
XU1355 n1449 n1450 VDD VSS INV_X32 
XU1356 n393 n1451 VDD VSS INV_X1 
XU1357 n1451 n1452 VDD VSS INV_X32 
XU1358 n1452 n1453 VDD VSS INV_X1 
XU1359 n1453 n1454 VDD VSS INV_X32 
XU1360 n1458 n1455 VDD VSS CLKBUF_X1 
XU1361 n1455 n1456 VDD VSS INV_X32 
XU1362 n1456 n1457 VDD VSS INV_X1 
XU1363 n380 n1458 VDD VSS INV_X1 
XU1364 n1457 n1459 VDD VSS INV_X32 
XU1365 n1465 n1460 VDD VSS INV_X1 
XU1366 n1460 n1461 VDD VSS INV_X32 
XU1367 n1464 n1462 VDD VSS INV_X32 
XU1368 n1462 n1463 VDD VSS INV_X1 
XU1369 n425 n1464 VDD VSS INV_X1 
XU1370 n1463 n1465 VDD VSS INV_X32 
XU1371 n652 n1466 VDD VSS INV_X32 
XU1372 n1466 n1467 VDD VSS INV_X1 
XU1373 n412 n1468 VDD VSS INV_X1 
XU1374 n1467 n1469 VDD VSS INV_X32 
XU1375 n163 n1470 VDD VSS CLKBUF_X1 
XU1376 n1474 n1471 VDD VSS CLKBUF_X1 
XU1377 n1471 n1472 VDD VSS INV_X32 
XU1378 n1472 n1473 VDD VSS INV_X1 
XU1379 n399 n1474 VDD VSS INV_X1 
XU1380 n1473 n1475 VDD VSS INV_X32 
XU1381 n1477 n1476 VDD VSS CLKBUF_X1 
XU1382 n386 n1477 VDD VSS INV_X1 
XU1383 n1476 n1478 VDD VSS INV_X32 
XU1384 n1478 n1479 VDD VSS INV_X1 
XU1385 n1479 n1480 VDD VSS INV_X32 
XU1386 n1486 n1481 VDD VSS INV_X1 
XU1387 n1481 n1482 VDD VSS INV_X32 
XU1388 n431 n1483 VDD VSS INV_X1 
XU1389 n1483 n1484 VDD VSS INV_X32 
XU1390 n1484 n1485 VDD VSS INV_X1 
XU1391 n1485 n1486 VDD VSS INV_X32 
XU1392 n1490 n1487 VDD VSS INV_X1 
XU1393 n1487 n1488 VDD VSS INV_X32 
XU1394 n418 n1489 VDD VSS INV_X1 
XU1395 n1489 n1490 VDD VSS INV_X32 
XU1396 n169 n1491 VDD VSS BUF_X1 
XU1397 n1493 n1492 VDD VSS CLKBUF_X1 
XU1398 n405 n1493 VDD VSS INV_X1 
XU1399 n1492 n1494 VDD VSS INV_X32 
XU1400 n1494 n1495 VDD VSS INV_X1 
XU1401 n1495 n1496 VDD VSS INV_X32 
XU1402 n1500 n1497 VDD VSS CLKBUF_X1 
XU1403 n392 n1498 VDD VSS INV_X1 
XU1404 n1498 n1499 VDD VSS INV_X32 
XU1405 n1499 n1500 VDD VSS INV_X1 
XU1406 n1497 n1501 VDD VSS INV_X32 
XU1407 n1505 n1502 VDD VSS CLKBUF_X1 
XU1408 n1502 n1503 VDD VSS INV_X32 
XU1409 n1503 n1504 VDD VSS INV_X1 
XU1410 n379 n1505 VDD VSS INV_X1 
XU1411 n1504 n1506 VDD VSS INV_X32 
XU1412 n1510 n1507 VDD VSS CLKBUF_X1 
XU1413 n1507 n1508 VDD VSS INV_X32 
XU1414 n1508 n1509 VDD VSS INV_X1 
XU1415 n424 n1510 VDD VSS INV_X1 
XU1416 n1509 n1511 VDD VSS INV_X32 
XU1417 n1513 n1512 VDD VSS CLKBUF_X1 
XU1418 n411 n1513 VDD VSS INV_X1 
XU1419 n1512 n1514 VDD VSS INV_X32 
XU1420 n1514 n1515 VDD VSS INV_X1 
XU1421 n1515 n1516 VDD VSS INV_X32 
XU1422 n1520 n1517 VDD VSS CLKBUF_X1 
XU1423 n1517 n1518 VDD VSS INV_X32 
XU1424 n1518 n1519 VDD VSS INV_X1 
XU1425 n398 n1520 VDD VSS INV_X1 
XU1426 n1519 n1521 VDD VSS INV_X32 
XU1427 n1525 n1522 VDD VSS CLKBUF_X1 
XU1428 n1522 n1523 VDD VSS INV_X32 
XU1429 n1523 n1524 VDD VSS INV_X1 
XU1430 n385 n1525 VDD VSS INV_X1 
XU1431 n1524 n1526 VDD VSS INV_X32 
XU1432 n1530 n1527 VDD VSS CLKBUF_X1 
XU1433 n1527 n1528 VDD VSS INV_X32 
XU1434 n1528 n1529 VDD VSS INV_X1 
XU1435 n430 n1530 VDD VSS INV_X1 
XU1436 n1529 n1531 VDD VSS INV_X32 
XU1437 n417 n1532 VDD VSS INV_X1 
XU1438 n1532 n1533 VDD VSS INV_X32 
XU1439 n1533 n1534 VDD VSS INV_X1 
XU1440 n1534 n1535 VDD VSS INV_X32 
XU1441 n168 n1536 VDD VSS INV_X1 
XU1442 n1536 n1537 VDD VSS INV_X32 
XU1443 n1539 n1538 VDD VSS CLKBUF_X1 
XU1444 n404 n1539 VDD VSS INV_X1 
XU1445 n1538 n1540 VDD VSS INV_X32 
XU1446 n1540 n1541 VDD VSS INV_X1 
XU1447 n1541 n1542 VDD VSS INV_X32 
XU1448 n1546 n1543 VDD VSS CLKBUF_X1 
XU1449 n391 n1544 VDD VSS INV_X1 
XU1450 n1544 n1545 VDD VSS INV_X32 
XU1451 n1545 n1546 VDD VSS INV_X1 
XU1452 n1543 n1547 VDD VSS INV_X32 
XU1453 n1551 n1548 VDD VSS CLKBUF_X1 
XU1454 n1548 n1549 VDD VSS INV_X32 
XU1455 n1549 n1550 VDD VSS INV_X1 
XU1456 n378 n1551 VDD VSS INV_X1 
XU1457 n1550 n1552 VDD VSS INV_X32 
XU1458 n1558 n1553 VDD VSS INV_X1 
XU1459 n1553 n1554 VDD VSS INV_X32 
XU1460 n1557 n1555 VDD VSS INV_X32 
XU1461 n1555 n1556 VDD VSS INV_X1 
XU1462 n423 n1557 VDD VSS INV_X1 
XU1463 n1556 n1558 VDD VSS INV_X32 
XU1464 n1564 n1559 VDD VSS INV_X1 
XU1465 n1559 n1560 VDD VSS INV_X32 
XU1466 n410 n1561 VDD VSS INV_X1 
XU1467 n1561 n1562 VDD VSS INV_X32 
XU1468 n1562 n1563 VDD VSS INV_X1 
XU1469 n1563 n1564 VDD VSS INV_X32 
XU1470 n1569 n1565 VDD VSS BUF_X1 
XU1471 n1568 n1566 VDD VSS INV_X32 
XU1472 n1566 n1567 VDD VSS INV_X1 
XU1473 n397 n1568 VDD VSS INV_X1 
XU1474 n1567 n1569 VDD VSS INV_X32 
XU1475 n673 n1570 VDD VSS INV_X32 
XU1476 n1570 n1571 VDD VSS INV_X1 
XU1477 n1572 n1573 VDD VSS INV_X1 
XU1478 n384 n1574 VDD VSS INV_X1 
XU1479 n1571 n1575 VDD VSS INV_X32 
XU1480 n1579 n1576 VDD VSS INV_X1 
XU1481 n1576 n1577 VDD VSS INV_X32 
XU1482 n429 n1578 VDD VSS INV_X1 
XU1483 n1578 n1579 VDD VSS INV_X32 
XU1484 n180 n1580 VDD VSS INV_X32 
XU1485 n1580 n1581 VDD VSS INV_X1 
XU1486 n1586 n1582 VDD VSS INV_X32 
XU1487 n1582 n1583 VDD VSS INV_X1 
XU1488 n1583 n1584 VDD VSS INV_X32 
XU1489 n1584 n1585 VDD VSS INV_X1 
XU1490 n416 n1586 VDD VSS INV_X1 
XU1491 n1585 n1587 VDD VSS INV_X32 
XU1492 n1589 n1588 VDD VSS CLKBUF_X1 
XU1493 n403 n1589 VDD VSS INV_X1 
XU1494 n1588 n1590 VDD VSS INV_X32 
XU1495 n1590 n1591 VDD VSS INV_X1 
XU1496 n1591 n1592 VDD VSS INV_X32 
XU1497 n1596 n1593 VDD VSS CLKBUF_X1 
XU1498 n1593 n1594 VDD VSS INV_X32 
XU1499 n1594 n1595 VDD VSS INV_X1 
XU1500 n390 n1596 VDD VSS INV_X1 
XU1501 n1595 n1597 VDD VSS INV_X32 
XU1502 n1601 n1598 VDD VSS CLKBUF_X1 
XU1503 n1598 n1599 VDD VSS INV_X32 
XU1504 n1599 n1600 VDD VSS INV_X1 
XU1505 n377 n1601 VDD VSS INV_X1 
XU1506 n1600 n1602 VDD VSS INV_X32 
XU1507 n1608 n1603 VDD VSS INV_X1 
XU1508 n1603 n1604 VDD VSS INV_X32 
XU1509 n1607 n1605 VDD VSS INV_X32 
XU1510 n1605 n1606 VDD VSS INV_X1 
XU1511 n422 n1607 VDD VSS INV_X1 
XU1512 n1606 n1608 VDD VSS INV_X32 
XU1513 n1610 n1609 VDD VSS CLKBUF_X1 
XU1514 n1613 n1610 VDD VSS INV_X1 
XU1515 n1609 n1611 VDD VSS INV_X32 
XU1516 n409 n1612 VDD VSS INV_X1 
XU1517 n1612 n1613 VDD VSS INV_X32 
XU1518 n1617 n1614 VDD VSS CLKBUF_X1 
XU1519 n1614 n1615 VDD VSS INV_X32 
XU1520 n1615 n1616 VDD VSS INV_X1 
XU1521 n396 n1617 VDD VSS INV_X1 
XU1522 n1616 n1618 VDD VSS INV_X32 
XU1523 n1622 n1619 VDD VSS CLKBUF_X1 
XU1524 n383 n1620 VDD VSS INV_X1 
XU1525 n1620 n1621 VDD VSS INV_X32 
XU1526 n1621 n1622 VDD VSS INV_X1 
XU1527 n1619 n1623 VDD VSS INV_X32 
XU1528 n1629 n1624 VDD VSS INV_X1 
XU1529 n1624 n1625 VDD VSS INV_X32 
XU1530 n1628 n1626 VDD VSS INV_X32 
XU1531 n1626 n1627 VDD VSS INV_X1 
XU1532 n428 n1628 VDD VSS INV_X1 
XU1533 n1627 n1629 VDD VSS INV_X32 
XU1534 n1635 n1630 VDD VSS INV_X1 
XU1535 n1630 n1631 VDD VSS INV_X32 
XU1536 n1634 n1632 VDD VSS INV_X32 
XU1537 n1632 n1633 VDD VSS INV_X1 
XU1538 n415 n1634 VDD VSS INV_X1 
XU1539 n1633 n1635 VDD VSS INV_X32 
XU1540 n682 n1636 VDD VSS INV_X32 
XU1541 n1636 n1637 VDD VSS INV_X1 
XU1542 n551 n1638 VDD VSS INV_X1 
XU1543 n1637 n1639 VDD VSS INV_X32 
XU1544 n55 n1640 VDD VSS CLKBUF_X1 
XU1545 n1643 n1641 VDD VSS INV_X32 
XU1546 n1641 n1642 VDD VSS INV_X1 
XU1547 n544 n1643 VDD VSS INV_X1 
XU1548 n1642 n1644 VDD VSS INV_X32 
XU1549 n48 n1645 VDD VSS INV_X1 
XU1550 n1645 n1646 VDD VSS INV_X32 
XU1551 n1648 n1647 VDD VSS CLKBUF_X1 
XU1552 n537 n1648 VDD VSS INV_X1 
XU1553 n1647 n1649 VDD VSS INV_X32 
XU1554 n1649 n1650 VDD VSS INV_X1 
XU1555 n1650 n1651 VDD VSS INV_X32 
XU1556 n1655 n1652 VDD VSS CLKBUF_X1 
XU1557 n1652 n1653 VDD VSS INV_X32 
XU1558 n1653 n1654 VDD VSS INV_X1 
XU1559 n530 n1655 VDD VSS INV_X1 
XU1560 n1654 n1656 VDD VSS INV_X32 
XU1561 n1658 n1657 VDD VSS CLKBUF_X1 
XU1562 n523 n1658 VDD VSS INV_X1 
XU1563 n1657 n1659 VDD VSS INV_X32 
XU1564 n1659 n1660 VDD VSS INV_X1 
XU1565 n1660 n1661 VDD VSS INV_X32 
XU1566 n1663 n1662 VDD VSS CLKBUF_X1 
XU1567 n516 n1663 VDD VSS INV_X1 
XU1568 n1662 n1664 VDD VSS INV_X32 
XU1569 n1664 n1665 VDD VSS INV_X1 
XU1570 n1665 n1666 VDD VSS INV_X32 
XU1571 n1670 n1667 VDD VSS CLKBUF_X1 
XU1572 n1667 n1668 VDD VSS INV_X32 
XU1573 n1668 n1669 VDD VSS INV_X1 
XU1574 n509 n1670 VDD VSS INV_X1 
XU1575 n1669 n1671 VDD VSS INV_X32 
XU1576 n689 n1672 VDD VSS INV_X32 
XU1577 n1672 n1673 VDD VSS INV_X1 
XU1578 n502 n1674 VDD VSS INV_X1 
XU1579 n1673 n1675 VDD VSS INV_X32 
XU1580 n6 n1676 VDD VSS BUF_X1 
XU1581 n1680 n1677 VDD VSS INV_X1 
XU1582 n691 n1678 VDD VSS INV_X32 
XU1583 n547 n1679 VDD VSS INV_X1 
XU1584 n1679 n1680 VDD VSS INV_X32 
XU1585 n51 n1681 VDD VSS BUF_X1 
XU1586 n1683 n1682 VDD VSS CLKBUF_X1 
XU1587 n540 n1683 VDD VSS INV_X1 
XU1588 n1682 n1684 VDD VSS INV_X32 
XU1589 n1684 n1685 VDD VSS INV_X1 
XU1590 n1685 n1686 VDD VSS INV_X32 
XU1591 n1692 n1687 VDD VSS INV_X1 
XU1592 n1687 n1688 VDD VSS INV_X32 
XU1593 n1691 n1689 VDD VSS INV_X32 
XU1594 n1689 n1690 VDD VSS INV_X1 
XU1595 n533 n1691 VDD VSS INV_X1 
XU1596 n1690 n1692 VDD VSS INV_X32 
XU1597 n1694 n1693 VDD VSS CLKBUF_X1 
XU1598 n526 n1694 VDD VSS INV_X1 
XU1599 n1693 n1695 VDD VSS INV_X32 
XU1600 n1695 n1696 VDD VSS INV_X1 
XU1601 n1696 n1697 VDD VSS INV_X32 
XU1602 n1701 n1698 VDD VSS CLKBUF_X1 
XU1603 n519 n1699 VDD VSS INV_X1 
XU1604 n1699 n1700 VDD VSS INV_X32 
XU1605 n1700 n1701 VDD VSS INV_X1 
XU1606 n1698 n1702 VDD VSS INV_X32 
XU1607 n1708 n1703 VDD VSS INV_X1 
XU1608 n1703 n1704 VDD VSS INV_X32 
XU1609 n512 n1705 VDD VSS INV_X1 
XU1610 n1705 n1706 VDD VSS INV_X32 
XU1611 n1706 n1707 VDD VSS INV_X1 
XU1612 n1707 n1708 VDD VSS INV_X32 
XU1613 n1712 n1709 VDD VSS CLKBUF_X1 
XU1614 n505 n1710 VDD VSS INV_X1 
XU1615 n1710 n1711 VDD VSS INV_X32 
XU1616 n1711 n1712 VDD VSS INV_X1 
XU1617 n1709 n1713 VDD VSS INV_X32 
XU1618 n498 n1714 VDD VSS INV_X1 
XU1619 n1714 n1715 VDD VSS INV_X32 
XU1620 n1715 n1716 VDD VSS INV_X1 
XU1621 n696 n1717 VDD VSS INV_X32 
XU1622 n2 n1718 VDD VSS INV_X1 
XU1623 n1718 n1719 VDD VSS INV_X8 
XU1624 n1723 n1720 VDD VSS CLKBUF_X1 
XU1625 n1720 n1721 VDD VSS INV_X32 
XU1626 n1721 n1722 VDD VSS INV_X1 
XU1627 n550 n1723 VDD VSS INV_X1 
XU1628 n1722 n1724 VDD VSS INV_X32 
XU1629 n699 n1725 VDD VSS INV_X32 
XU1630 n1725 n1726 VDD VSS INV_X1 
XU1631 n543 n1727 VDD VSS INV_X1 
XU1632 n1726 n1728 VDD VSS INV_X32 
XU1633 n47 n1729 VDD VSS BUF_X1 
XU1634 n1735 n1730 VDD VSS INV_X1 
XU1635 n1730 n1731 VDD VSS INV_X32 
XU1636 n1734 n1732 VDD VSS INV_X32 
XU1637 n1732 n1733 VDD VSS INV_X1 
XU1638 n536 n1734 VDD VSS INV_X1 
XU1639 n1733 n1735 VDD VSS INV_X32 
XU1640 n1739 n1736 VDD VSS CLKBUF_X1 
XU1641 n1736 n1737 VDD VSS INV_X32 
XU1642 n1737 n1738 VDD VSS INV_X1 
XU1643 n529 n1739 VDD VSS INV_X1 
XU1644 n1738 n1740 VDD VSS INV_X32 
XU1645 n1744 n1741 VDD VSS CLKBUF_X1 
XU1646 n1741 n1742 VDD VSS INV_X32 
XU1647 n1742 n1743 VDD VSS INV_X1 
XU1648 n522 n1744 VDD VSS INV_X1 
XU1649 n1743 n1745 VDD VSS INV_X32 
XU1650 n1749 n1746 VDD VSS CLKBUF_X1 
XU1651 n1746 n1747 VDD VSS INV_X32 
XU1652 n1747 n1748 VDD VSS INV_X1 
XU1653 n515 n1749 VDD VSS INV_X1 
XU1654 n1748 n1750 VDD VSS INV_X32 
XU1655 n1754 n1751 VDD VSS CLKBUF_X1 
XU1656 n508 n1752 VDD VSS INV_X1 
XU1657 n1752 n1753 VDD VSS INV_X32 
XU1658 n1753 n1754 VDD VSS INV_X1 
XU1659 n1751 n1755 VDD VSS INV_X32 
XU1660 n1757 n1756 VDD VSS CLKBUF_X1 
XU1661 n501 n1757 VDD VSS INV_X1 
XU1662 n1756 n1758 VDD VSS INV_X32 
XU1663 n1758 n1759 VDD VSS INV_X1 
XU1664 n1759 n1760 VDD VSS INV_X32 
XU1665 n1764 n1761 VDD VSS INV_X1 
XU1666 n706 n1762 VDD VSS INV_X32 
XU1667 n546 n1763 VDD VSS INV_X1 
XU1668 n1763 n1764 VDD VSS INV_X32 
XU1669 n50 n1765 VDD VSS BUF_X1 
XU1670 n1767 n1766 VDD VSS CLKBUF_X1 
XU1671 n539 n1767 VDD VSS INV_X1 
XU1672 n1766 n1768 VDD VSS INV_X32 
XU1673 n1768 n1769 VDD VSS INV_X1 
XU1674 n1769 n1770 VDD VSS INV_X32 
XU1675 n1776 n1771 VDD VSS INV_X1 
XU1676 n1771 n1772 VDD VSS INV_X32 
XU1677 n1775 n1773 VDD VSS INV_X32 
XU1678 n1773 n1774 VDD VSS INV_X1 
XU1679 n532 n1775 VDD VSS INV_X1 
XU1680 n1774 n1776 VDD VSS INV_X32 
XU1681 n1780 n1777 VDD VSS CLKBUF_X1 
XU1682 n1777 n1778 VDD VSS INV_X32 
XU1683 n1778 n1779 VDD VSS INV_X1 
XU1684 n525 n1780 VDD VSS INV_X1 
XU1685 n1779 n1781 VDD VSS INV_X32 
XU1686 n1785 n1782 VDD VSS CLKBUF_X1 
XU1687 n518 n1783 VDD VSS INV_X1 
XU1688 n1783 n1784 VDD VSS INV_X32 
XU1689 n1784 n1785 VDD VSS INV_X1 
XU1690 n1782 n1786 VDD VSS INV_X32 
XU1691 n1791 n1787 VDD VSS BUF_X1 
XU1692 n1790 n1788 VDD VSS INV_X32 
XU1693 n1788 n1789 VDD VSS INV_X1 
XU1694 n511 n1790 VDD VSS INV_X1 
XU1695 n1789 n1791 VDD VSS INV_X32 
XU1696 n504 n1792 VDD VSS INV_X1 
XU1697 n1792 n1793 VDD VSS INV_X32 
XU1698 n1793 n1794 VDD VSS INV_X1 
XU1699 n1794 n1795 VDD VSS INV_X32 
XU1700 n15 n1796 VDD VSS INV_X32 
XU1701 n1796 n1797 VDD VSS INV_X1 
XU1702 n1801 n1798 VDD VSS CLKBUF_X1 
XU1703 n1798 n1799 VDD VSS INV_X32 
XU1704 n1799 n1800 VDD VSS INV_X1 
XU1705 n497 n1801 VDD VSS INV_X1 
XU1706 n1800 n1802 VDD VSS INV_X32 
XU1707 n1808 n1803 VDD VSS INV_X1 
XU1708 n1803 n1804 VDD VSS INV_X32 
XU1709 n1807 n1805 VDD VSS INV_X32 
XU1710 n1805 n1806 VDD VSS INV_X1 
XU1711 n549 n1807 VDD VSS INV_X1 
XU1712 n1806 n1808 VDD VSS INV_X32 
XU1713 n1810 n1809 VDD VSS CLKBUF_X1 
XU1714 n542 n1810 VDD VSS INV_X1 
XU1715 n1809 n1811 VDD VSS INV_X32 
XU1716 n1811 n1812 VDD VSS INV_X1 
XU1717 n1812 n1813 VDD VSS INV_X32 
XU1718 n1817 n1814 VDD VSS CLKBUF_X1 
XU1719 n1814 n1815 VDD VSS INV_X32 
XU1720 n1815 n1816 VDD VSS INV_X1 
XU1721 n535 n1817 VDD VSS INV_X1 
XU1722 n1816 n1818 VDD VSS INV_X32 
XU1723 n1822 n1819 VDD VSS CLKBUF_X1 
XU1724 n528 n1820 VDD VSS INV_X1 
XU1725 n1820 n1821 VDD VSS INV_X32 
XU1726 n1821 n1822 VDD VSS INV_X1 
XU1727 n1819 n1823 VDD VSS INV_X32 
XU1728 n1827 n1824 VDD VSS CLKBUF_X1 
XU1729 n1824 n1825 VDD VSS INV_X32 
XU1730 n1825 n1826 VDD VSS INV_X1 
XU1731 n521 n1827 VDD VSS INV_X1 
XU1732 n1826 n1828 VDD VSS INV_X32 
XU1733 n1832 n1829 VDD VSS CLKBUF_X1 
XU1734 n1829 n1830 VDD VSS INV_X32 
XU1735 n1830 n1831 VDD VSS INV_X1 
XU1736 n514 n1832 VDD VSS INV_X1 
XU1737 n1831 n1833 VDD VSS INV_X32 
XU1738 n1839 n1834 VDD VSS INV_X1 
XU1739 n1834 n1835 VDD VSS INV_X32 
XU1740 n507 n1836 VDD VSS INV_X1 
XU1741 n1836 n1837 VDD VSS INV_X32 
XU1742 n1837 n1838 VDD VSS INV_X1 
XU1743 n1838 n1839 VDD VSS INV_X32 
XU1744 n1843 n1840 VDD VSS CLKBUF_X1 
XU1745 n1840 n1841 VDD VSS INV_X32 
XU1746 n1841 n1842 VDD VSS INV_X1 
XU1747 n500 n1843 VDD VSS INV_X1 
XU1748 n1842 n1844 VDD VSS INV_X32 
XU1749 n1848 n1845 VDD VSS CLKBUF_X1 
XU1750 n1845 n1846 VDD VSS INV_X32 
XU1751 n1846 n1847 VDD VSS INV_X1 
XU1752 n545 n1848 VDD VSS INV_X1 
XU1753 n1847 n1849 VDD VSS INV_X32 
XU1754 n1851 n1850 VDD VSS CLKBUF_X1 
XU1755 n1854 n1851 VDD VSS INV_X1 
XU1756 n1850 n1852 VDD VSS INV_X32 
XU1757 n538 n1853 VDD VSS INV_X1 
XU1758 n1853 n1854 VDD VSS INV_X32 
XU1759 n1858 n1855 VDD VSS CLKBUF_X1 
XU1760 n531 n1856 VDD VSS INV_X1 
XU1761 n1856 n1857 VDD VSS INV_X32 
XU1762 n1857 n1858 VDD VSS INV_X1 
XU1763 n1855 n1859 VDD VSS INV_X32 
XU1764 n1865 n1860 VDD VSS INV_X1 
XU1765 n1860 n1861 VDD VSS INV_X32 
XU1766 n1864 n1862 VDD VSS INV_X32 
XU1767 n1862 n1863 VDD VSS INV_X1 
XU1768 n524 n1864 VDD VSS INV_X1 
XU1769 n1863 n1865 VDD VSS INV_X32 
XU1770 n1867 n1866 VDD VSS CLKBUF_X1 
XU1771 n1870 n1867 VDD VSS INV_X1 
XU1772 n1866 n1868 VDD VSS INV_X32 
XU1773 n517 n1869 VDD VSS INV_X1 
XU1774 n1869 n1870 VDD VSS INV_X32 
XU1775 n1874 n1871 VDD VSS CLKBUF_X1 
XU1776 n1871 n1872 VDD VSS INV_X32 
XU1777 n1872 n1873 VDD VSS INV_X1 
XU1778 n510 n1874 VDD VSS INV_X1 
XU1779 n1873 n1875 VDD VSS INV_X32 
XU1780 n503 n1876 VDD VSS INV_X1 
XU1781 n1876 n1877 VDD VSS INV_X32 
XU1782 n1877 n1878 VDD VSS INV_X1 
XU1783 n723 n1879 VDD VSS INV_X32 
XU1784 n7 n1880 VDD VSS INV_X1 
XU1785 n1880 n1881 VDD VSS INV_X8 
XU1786 n725 n1882 VDD VSS INV_X32 
XU1787 n1882 n1883 VDD VSS INV_X1 
XU1788 n548 n1884 VDD VSS INV_X1 
XU1789 n1883 n1885 VDD VSS INV_X32 
XU1790 n52 n1886 VDD VSS CLKBUF_X1 
XU1791 n1888 n1887 VDD VSS CLKBUF_X1 
XU1792 n541 n1888 VDD VSS INV_X1 
XU1793 n1887 n1889 VDD VSS INV_X32 
XU1794 n1889 n1890 VDD VSS INV_X1 
XU1795 n1890 n1891 VDD VSS INV_X32 
XU1796 n1895 n1892 VDD VSS CLKBUF_X1 
XU1797 n534 n1893 VDD VSS INV_X1 
XU1798 n1893 n1894 VDD VSS INV_X32 
XU1799 n1894 n1895 VDD VSS INV_X1 
XU1800 n1892 n1896 VDD VSS INV_X32 
XU1801 n1900 n1897 VDD VSS CLKBUF_X1 
XU1802 n527 n1898 VDD VSS INV_X1 
XU1803 n1898 n1899 VDD VSS INV_X32 
XU1804 n1899 n1900 VDD VSS INV_X1 
XU1805 n1897 n1901 VDD VSS INV_X32 
XU1806 n1903 n1902 VDD VSS CLKBUF_X1 
XU1807 n1906 n1903 VDD VSS INV_X1 
XU1808 n1902 n1904 VDD VSS INV_X32 
XU1809 n520 n1905 VDD VSS INV_X1 
XU1810 n1905 n1906 VDD VSS INV_X32 
XU1811 n1908 n1907 VDD VSS CLKBUF_X1 
XU1812 n513 n1908 VDD VSS INV_X1 
XU1813 n1907 n1909 VDD VSS INV_X32 
XU1814 n1909 n1910 VDD VSS INV_X1 
XU1815 n1910 n1911 VDD VSS INV_X32 
XU1816 n1915 n1912 VDD VSS CLKBUF_X1 
XU1817 n1912 n1913 VDD VSS INV_X32 
XU1818 n1913 n1914 VDD VSS INV_X1 
XU1819 n506 n1915 VDD VSS INV_X1 
XU1820 n1914 n1916 VDD VSS INV_X32 
XU1821 n1920 n1917 VDD VSS CLKBUF_X1 
XU1822 n1917 n1918 VDD VSS INV_X32 
XU1823 n1918 n1919 VDD VSS INV_X1 
XU1824 n499 n1920 VDD VSS INV_X1 
XU1825 n1919 n1921 VDD VSS INV_X32 
XU1826 n1925 n1922 VDD VSS CLKBUF_X1 
XU1827 n1922 n1923 VDD VSS INV_X32 
XU1828 n1923 n1924 VDD VSS INV_X1 
XU1829 n496 n1925 VDD VSS INV_X1 
XU1830 n1924 n1926 VDD VSS INV_X32 
XU1831 n736 n1927 VDD VSS INV_X32 
XU1832 n1927 n1928 VDD VSS INV_X1 
XU1833 n472 n1929 VDD VSS INV_X1 
XU1834 n1928 n1930 VDD VSS INV_X32 
XU1835 n99 n1931 VDD VSS BUF_X1 
XU1836 n1937 n1932 VDD VSS INV_X1 
XU1837 n1932 n1933 VDD VSS INV_X32 
XU1838 n448 n1934 VDD VSS INV_X1 
XU1839 n1934 n1935 VDD VSS INV_X32 
XU1840 n1935 n1936 VDD VSS INV_X1 
XU1841 n1936 n1937 VDD VSS INV_X32 
XU1842 n1941 n1938 VDD VSS CLKBUF_X1 
XU1843 n482 n1939 VDD VSS INV_X1 
XU1844 n1939 n1940 VDD VSS INV_X32 
XU1845 n1940 n1941 VDD VSS INV_X1 
XU1846 n1938 n1942 VDD VSS INV_X32 
XU1847 n1946 n1943 VDD VSS CLKBUF_X1 
XU1848 n1943 n1944 VDD VSS INV_X32 
XU1849 n1944 n1945 VDD VSS INV_X1 
XU1850 n458 n1946 VDD VSS INV_X1 
XU1851 n1945 n1947 VDD VSS INV_X32 
XU1852 n1953 n1948 VDD VSS INV_X1 
XU1853 n1948 n1949 VDD VSS INV_X32 
XU1854 n1952 n1950 VDD VSS INV_X32 
XU1855 n1950 n1951 VDD VSS INV_X1 
XU1856 n434 n1952 VDD VSS INV_X1 
XU1857 n1951 n1953 VDD VSS INV_X32 
XU1858 n1957 n1954 VDD VSS CLKBUF_X1 
XU1859 n1954 n1955 VDD VSS INV_X32 
XU1860 n1955 n1956 VDD VSS INV_X1 
XU1861 n492 n1957 VDD VSS INV_X1 
XU1862 n1956 n1958 VDD VSS INV_X32 
XU1863 n1962 n1959 VDD VSS CLKBUF_X1 
XU1864 n1959 n1960 VDD VSS INV_X32 
XU1865 n1960 n1961 VDD VSS INV_X1 
XU1866 n468 n1962 VDD VSS INV_X1 
XU1867 n1961 n1963 VDD VSS INV_X32 
XU1868 n1967 n1964 VDD VSS CLKBUF_X1 
XU1869 n444 n1965 VDD VSS INV_X1 
XU1870 n1965 n1966 VDD VSS INV_X32 
XU1871 n1966 n1967 VDD VSS INV_X1 
XU1872 n1964 n1968 VDD VSS INV_X32 
XU1873 n478 n1969 VDD VSS INV_X1 
XU1874 n1969 n1970 VDD VSS INV_X32 
XU1875 n1970 n1971 VDD VSS INV_X1 
XU1876 n1971 n1972 VDD VSS INV_X32 
XU1877 n1973 n1974 VDD VSS INV_X1 
XU1878 n1980 n1975 VDD VSS INV_X1 
XU1879 n1975 n1976 VDD VSS INV_X32 
XU1880 n1979 n1977 VDD VSS INV_X32 
XU1881 n1977 n1978 VDD VSS INV_X1 
XU1882 n454 n1979 VDD VSS INV_X1 
XU1883 n1978 n1980 VDD VSS INV_X32 
XU1884 n1984 n1981 VDD VSS CLKBUF_X1 
XU1885 n1981 n1982 VDD VSS INV_X32 
XU1886 n1982 n1983 VDD VSS INV_X1 
XU1887 n493 n1984 VDD VSS INV_X1 
XU1888 n1983 n1985 VDD VSS INV_X32 
XU1889 n1987 n1986 VDD VSS CLKBUF_X1 
XU1890 n469 n1987 VDD VSS INV_X1 
XU1891 n1986 n1988 VDD VSS INV_X32 
XU1892 n1988 n1989 VDD VSS INV_X1 
XU1893 n1989 n1990 VDD VSS INV_X32 
XU1894 n1994 n1991 VDD VSS CLKBUF_X1 
XU1895 n1991 n1992 VDD VSS INV_X32 
XU1896 n1992 n1993 VDD VSS INV_X1 
XU1897 n445 n1994 VDD VSS INV_X1 
XU1898 n1993 n1995 VDD VSS INV_X32 
XU1899 n1999 n1996 VDD VSS INV_X1 
XU1900 n1996 n1997 VDD VSS INV_X32 
XU1901 n479 n1998 VDD VSS INV_X1 
XU1902 n1998 n1999 VDD VSS INV_X32 
XU1903 n106 n2000 VDD VSS INV_X32 
XU1904 n2000 n2001 VDD VSS INV_X1 
XU1905 n2005 n2002 VDD VSS INV_X32 
XU1906 n2002 n2003 VDD VSS INV_X1 
XU1907 n2006 n2004 VDD VSS INV_X32 
XU1908 n2004 n2005 VDD VSS INV_X1 
XU1909 n455 n2006 VDD VSS INV_X1 
XU1910 n2003 n2007 VDD VSS INV_X32 
XU1911 n2011 n2008 VDD VSS CLKBUF_X1 
XU1912 n2008 n2009 VDD VSS INV_X32 
XU1913 n2009 n2010 VDD VSS INV_X1 
XU1914 n494 n2011 VDD VSS INV_X1 
XU1915 n2010 n2012 VDD VSS INV_X32 
XU1916 n2025 n2013 VDD VSS CLKBUF_X1 
XU1917 n2015 n2014 VDD VSS CLKBUF_X1 
XU1918 n2013 n2015 VDD VSS INV_X32 
XU1919 n2014 data_out[0] VDD VSS INV_X32 
XU1920 n2026 n2017 VDD VSS CLKBUF_X1 
XU1921 n2017 n2018 VDD VSS INV_X32 
XU1922 n2018 data_out[6] VDD VSS INV_X1 
XU1923 n2024 n2020 VDD VSS CLKBUF_X1 
XU1924 n2022 n2021 VDD VSS CLKBUF_X1 
XU1925 n2020 n2022 VDD VSS INV_X32 
XU1926 n2021 data_out[14] VDD VSS INV_X32 
XU722 n811 n812 VDD VSS INV_X2 
XU1927 n812 n2027 VDD VSS BUF_X1 
XU1928 n1071 n2028 VDD VSS BUF_X1 
XU1929 n830 n2029 VDD VSS BUF_X1 
XU1930 n1045 n2030 VDD VSS BUF_X1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW01_add_1 CI CO VDD VSS SUM[31] SUM[30] SUM[29] SUM[28] 
+ SUM[27] SUM[26] SUM[25] SUM[24] SUM[23] SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] 
+ SUM[17] SUM[16] SUM[15] SUM[14] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] 
+ B[23] B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] 
+ B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[31] A[30] A[29] A[28] 
+ A[27] A[26] A[25] A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] 
+ A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU7 n30 n3 VDD VSS INV_X1 
XU6 n38 n5 VDD VSS INV_X1 
XU5 n46 n7 VDD VSS INV_X1 
XU4 n54 n9 VDD VSS INV_X1 
XU3 n62 n11 VDD VSS INV_X1 
XU2 n70 n13 VDD VSS INV_X1 
XU100 B[15] A[15] n80 VDD VSS NOR2_X1 
XU99 B[15] A[15] n82 VDD VSS NAND2_X1 
XU98 n16 n82 n83 VDD VSS NAND2_X1 
XU97 n81 n83 n155 VDD VSS XOR2_X1 
XU96 n82 n80 n81 n76 VDD VSS OAI21_X1 
XU95 B[16] A[16] n77 VDD VSS AND2_X1 
XU94 B[16] A[16] n78 VDD VSS NOR2_X1 
XU93 n77 n78 n79 VDD VSS NOR2_X1 
XU92 n76 n79 n147 VDD VSS XOR2_X1 
XU91 B[17] A[17] n72 VDD VSS NOR2_X1 
XU90 B[17] A[17] n74 VDD VSS NAND2_X1 
XU89 n14 n74 n75 VDD VSS NAND2_X1 
XU88 n77 n15 n76 n73 VDD VSS AOI21_X1 
XU87 n75 n73 n148 VDD VSS XOR2_X1 
XU86 n74 n72 n73 n68 VDD VSS OAI21_X1 
XU85 B[18] A[18] n69 VDD VSS AND2_X1 
XU84 B[18] A[18] n70 VDD VSS NOR2_X1 
XU83 n69 n70 n71 VDD VSS NOR2_X1 
XU82 n68 n71 n149 VDD VSS XOR2_X1 
XU81 B[19] A[19] n64 VDD VSS NOR2_X1 
XU80 B[19] A[19] n66 VDD VSS NAND2_X1 
XU79 n12 n66 n67 VDD VSS NAND2_X1 
XU78 n69 n13 n68 n65 VDD VSS AOI21_X1 
XU77 n67 n65 n150 VDD VSS XOR2_X1 
XU76 n66 n64 n65 n60 VDD VSS OAI21_X1 
XU75 B[20] A[20] n61 VDD VSS AND2_X1 
XU74 B[20] A[20] n62 VDD VSS NOR2_X1 
XU73 n61 n62 n63 VDD VSS NOR2_X1 
XU72 n60 n63 n151 VDD VSS XOR2_X1 
XU71 B[21] A[21] n56 VDD VSS NOR2_X1 
XU70 B[21] A[21] n58 VDD VSS NAND2_X1 
XU69 n10 n58 n59 VDD VSS NAND2_X1 
XU68 n61 n11 n60 n57 VDD VSS AOI21_X1 
XU67 n59 n57 n152 VDD VSS XOR2_X1 
XU66 n58 n56 n57 n52 VDD VSS OAI21_X1 
XU65 B[22] A[22] n53 VDD VSS AND2_X1 
XU64 B[22] A[22] n54 VDD VSS NOR2_X1 
XU63 n53 n54 n55 VDD VSS NOR2_X1 
XU62 n52 n55 n153 VDD VSS XOR2_X1 
XU61 B[23] A[23] n48 VDD VSS NOR2_X1 
XU60 B[23] A[23] n50 VDD VSS NAND2_X1 
XU59 n8 n85 n51 VDD VSS NAND2_X1 
XU58 n53 n9 n52 n49 VDD VSS AOI21_X1 
XU57 n51 n49 n154 VDD VSS XOR2_X1 
XU56 n85 n48 n49 n44 VDD VSS OAI21_X1 
XU55 B[24] A[24] n45 VDD VSS AND2_X1 
XU54 B[24] A[24] n46 VDD VSS NOR2_X1 
XU53 n45 n46 n47 VDD VSS NOR2_X1 
XU52 n44 n47 n139 VDD VSS XOR2_X1 
XU51 B[25] A[25] n40 VDD VSS NOR2_X1 
XU50 B[25] A[25] n42 VDD VSS NAND2_X1 
XU49 n6 n42 n43 VDD VSS NAND2_X1 
XU48 n45 n7 n44 n41 VDD VSS AOI21_X1 
XU47 n43 n41 n140 VDD VSS XOR2_X1 
XU46 n42 n40 n41 n36 VDD VSS OAI21_X1 
XU45 B[26] A[26] n37 VDD VSS AND2_X1 
XU44 B[26] A[26] n38 VDD VSS NOR2_X1 
XU43 n37 n38 n39 VDD VSS NOR2_X1 
XU42 n36 n39 n141 VDD VSS XOR2_X1 
XU41 B[27] A[27] n32 VDD VSS NOR2_X1 
XU40 B[27] A[27] n34 VDD VSS NAND2_X1 
XU39 n4 n34 n35 VDD VSS NAND2_X1 
XU38 n37 n5 n36 n33 VDD VSS AOI21_X1 
XU37 n35 n33 n142 VDD VSS XOR2_X1 
XU36 n34 n32 n33 n28 VDD VSS OAI21_X1 
XU35 B[28] A[28] n29 VDD VSS AND2_X1 
XU34 B[28] A[28] n30 VDD VSS NOR2_X1 
XU33 n29 n30 n31 VDD VSS NOR2_X1 
XU32 n28 n31 n143 VDD VSS XOR2_X1 
XU31 B[29] A[29] n24 VDD VSS NOR2_X1 
XU30 B[29] A[29] n26 VDD VSS NAND2_X1 
XU29 n2 n26 n27 VDD VSS NAND2_X1 
XU28 n29 n3 n28 n25 VDD VSS AOI21_X1 
XU27 n27 n25 n144 VDD VSS XOR2_X1 
XU26 n26 n24 n25 n20 VDD VSS OAI21_X1 
XU25 B[30] A[30] n21 VDD VSS AND2_X1 
XU24 B[30] A[30] n22 VDD VSS NOR2_X1 
XU23 n21 n22 n23 VDD VSS NOR2_X1 
XU22 n20 n23 n145 VDD VSS XOR2_X1 
XU21 B[31] A[31] n18 VDD VSS XNOR2_X1 
XU20 n21 n20 n1 n19 VDD VSS AOI21_X1 
XU19 n18 n19 n146 VDD VSS XOR2_X1 
XU18 n126 SUM[14] VDD VSS INV_X1 
XU17 n80 n16 VDD VSS INV_X1 
XU16 n78 n15 VDD VSS INV_X1 
XU15 n22 n1 VDD VSS INV_X1 
XU14 n40 n6 VDD VSS INV_X1 
XU13 n48 n8 VDD VSS INV_X1 
XU12 n56 n10 VDD VSS INV_X1 
XU11 n64 n12 VDD VSS INV_X1 
XU10 n72 n14 VDD VSS INV_X1 
XU9 n24 n2 VDD VSS INV_X1 
XU8 n32 n4 VDD VSS INV_X1 
XU102 B[14] A[14] n81 VDD VSS NAND2_X1 
XU101 n81 B[14] A[14] n84 VDD VSS OAI21_X1 
XU1 n91 SUM[26] VDD VSS BUF_X1 
XU103 n50 n85 VDD VSS BUF_X1 
XU104 n107 SUM[20] VDD VSS BUF_X1 
XU105 n143 n137 VDD VSS INV_X2 
XU106 n145 n131 VDD VSS INV_X4 
XU107 n144 n134 VDD VSS INV_X4 
XU108 n153 n102 VDD VSS INV_X1 
XU109 n154 n99 VDD VSS INV_X1 
XU110 n89 n87 VDD VSS INV_X1 
XU111 n87 SUM[27] VDD VSS INV_X8 
XU112 n142 n89 VDD VSS BUF_X32 
XU113 n92 n90 VDD VSS INV_X1 
XU114 n90 n91 VDD VSS INV_X4 
XU115 n141 n92 VDD VSS BUF_X32 
XU116 n95 n93 VDD VSS INV_X1 
XU117 n93 SUM[25] VDD VSS INV_X8 
XU118 n140 n95 VDD VSS BUF_X32 
XU119 n97 SUM[24] VDD VSS BUF_X1 
XU120 n139 n97 VDD VSS BUF_X32 
XU121 n100 SUM[23] VDD VSS BUF_X1 
XU122 n99 n100 VDD VSS INV_X32 
XU123 n103 SUM[22] VDD VSS BUF_X1 
XU124 n102 n103 VDD VSS INV_X32 
XU125 n106 n104 VDD VSS INV_X1 
XU126 n104 SUM[21] VDD VSS INV_X8 
XU127 n152 n106 VDD VSS BUF_X32 
XU128 n108 n107 VDD VSS CLKBUF_X1 
XU129 n151 n108 VDD VSS BUF_X32 
XU130 n111 n109 VDD VSS INV_X1 
XU131 n109 SUM[19] VDD VSS INV_X8 
XU132 n150 n111 VDD VSS BUF_X32 
XU133 n114 n112 VDD VSS INV_X1 
XU134 n112 SUM[18] VDD VSS INV_X8 
XU135 n149 n114 VDD VSS BUF_X32 
XU136 n117 n115 VDD VSS INV_X1 
XU137 n115 SUM[17] VDD VSS INV_X8 
XU138 n148 n117 VDD VSS BUF_X32 
XU139 n120 SUM[16] VDD VSS BUF_X1 
XU140 n147 n119 VDD VSS INV_X1 
XU141 n119 n120 VDD VSS INV_X32 
XU142 n123 SUM[15] VDD VSS BUF_X1 
XU143 n155 n122 VDD VSS INV_X1 
XU144 n122 n123 VDD VSS INV_X32 
XU145 n125 n124 VDD VSS CLKBUF_X1 
XU146 n84 n125 VDD VSS INV_X1 
XU147 n124 n126 VDD VSS INV_X32 
XU148 n128 n127 VDD VSS CLKBUF_X1 
XU149 n146 n128 VDD VSS INV_X1 
XU150 n127 SUM[31] VDD VSS INV_X32 
XU151 n131 n130 VDD VSS BUF_X1 
XU152 n130 SUM[30] VDD VSS INV_X32 
XU153 n134 n133 VDD VSS BUF_X1 
XU154 n133 SUM[29] VDD VSS INV_X32 
XU155 n137 n136 VDD VSS BUF_X1 
XU156 n136 SUM[28] VDD VSS INV_X32 
.ENDS

.SUBCKT gng_smul_16_18_DW01_add_0 CI CO VDD VSS SUM[31] SUM[30] SUM[29] SUM[28] SUM[27] 
+ SUM[26] SUM[25] SUM[24] SUM[23] SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] SUM[17] 
+ SUM[16] SUM[15] SUM[14] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] B[23] 
+ B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] 
+ B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[31] A[30] A[29] A[28] A[27] 
+ A[26] A[25] A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] 
+ A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU44 B[26] A[26] n38 VDD VSS NOR2_X1 
XU43 n37 n38 n39 VDD VSS NOR2_X1 
XU42 n36 n39 n129 VDD VSS XOR2_X1 
XU41 B[27] A[27] n32 VDD VSS NOR2_X1 
XU40 B[27] A[27] n34 VDD VSS NAND2_X1 
XU39 n4 n34 n35 VDD VSS NAND2_X1 
XU38 n37 n5 n36 n33 VDD VSS AOI21_X1 
XU37 n35 n33 n130 VDD VSS XOR2_X1 
XU36 n34 n32 n33 n28 VDD VSS OAI21_X1 
XU35 B[28] A[28] n29 VDD VSS AND2_X1 
XU34 B[28] A[28] n30 VDD VSS NOR2_X1 
XU33 n29 n30 n31 VDD VSS NOR2_X1 
XU32 n28 n31 n131 VDD VSS XOR2_X1 
XU31 B[29] A[29] n24 VDD VSS NOR2_X1 
XU30 B[29] A[29] n26 VDD VSS NAND2_X1 
XU29 n2 n26 n27 VDD VSS NAND2_X1 
XU28 n29 n3 n28 n25 VDD VSS AOI21_X1 
XU27 n27 n25 n132 VDD VSS XOR2_X1 
XU26 n26 n24 n25 n20 VDD VSS OAI21_X1 
XU25 B[30] A[30] n21 VDD VSS AND2_X1 
XU24 B[30] A[30] n22 VDD VSS NOR2_X1 
XU23 n21 n22 n23 VDD VSS NOR2_X1 
XU22 n20 n23 n133 VDD VSS XOR2_X1 
XU21 B[31] A[31] n18 VDD VSS XNOR2_X1 
XU20 n21 n20 n1 n19 VDD VSS AOI21_X1 
XU19 n18 n19 SUM[31] VDD VSS XOR2_X1 
XU18 n84 SUM[14] VDD VSS INV_X1 
XU17 n80 n16 VDD VSS INV_X1 
XU16 n78 n15 VDD VSS INV_X1 
XU15 n22 n1 VDD VSS INV_X1 
XU14 n40 n6 VDD VSS INV_X1 
XU13 n48 n8 VDD VSS INV_X1 
XU12 n56 n10 VDD VSS INV_X1 
XU11 n64 n12 VDD VSS INV_X1 
XU10 n72 n14 VDD VSS INV_X1 
XU9 n24 n2 VDD VSS INV_X1 
XU8 n32 n4 VDD VSS INV_X1 
XU7 n30 n3 VDD VSS INV_X1 
XU6 n38 n5 VDD VSS INV_X1 
XU5 n46 n7 VDD VSS INV_X1 
XU4 n54 n9 VDD VSS INV_X1 
XU3 n62 n11 VDD VSS INV_X1 
XU2 n70 n13 VDD VSS INV_X1 
XU102 B[14] A[14] n81 VDD VSS NAND2_X1 
XU101 n81 B[14] A[14] n84 VDD VSS OAI21_X1 
XU100 B[15] A[15] n80 VDD VSS NOR2_X1 
XU99 B[15] A[15] n82 VDD VSS NAND2_X1 
XU98 n16 n82 n83 VDD VSS NAND2_X1 
XU97 n81 n83 SUM[15] VDD VSS XOR2_X1 
XU96 n82 n80 n81 n76 VDD VSS OAI21_X1 
XU95 B[16] A[16] n77 VDD VSS AND2_X1 
XU94 B[16] A[16] n78 VDD VSS NOR2_X1 
XU93 n77 n78 n79 VDD VSS NOR2_X1 
XU92 n76 n79 SUM[16] VDD VSS XOR2_X1 
XU91 B[17] A[17] n72 VDD VSS NOR2_X1 
XU90 B[17] A[17] n74 VDD VSS NAND2_X1 
XU89 n14 n74 n75 VDD VSS NAND2_X1 
XU88 n77 n15 n76 n73 VDD VSS AOI21_X1 
XU87 n75 n73 n134 VDD VSS XOR2_X1 
XU86 n74 n72 n73 n68 VDD VSS OAI21_X1 
XU85 B[18] A[18] n69 VDD VSS AND2_X1 
XU84 B[18] A[18] n70 VDD VSS NOR2_X1 
XU83 n69 n70 n71 VDD VSS NOR2_X1 
XU82 n68 n71 n135 VDD VSS XOR2_X1 
XU81 B[19] A[19] n64 VDD VSS NOR2_X1 
XU80 B[19] A[19] n66 VDD VSS NAND2_X1 
XU79 n12 n66 n67 VDD VSS NAND2_X1 
XU78 n69 n13 n68 n65 VDD VSS AOI21_X1 
XU77 n67 n65 n136 VDD VSS XOR2_X1 
XU76 n66 n64 n65 n60 VDD VSS OAI21_X1 
XU75 B[20] A[20] n61 VDD VSS AND2_X1 
XU74 B[20] A[20] n62 VDD VSS NOR2_X1 
XU73 n61 n62 n63 VDD VSS NOR2_X1 
XU72 n60 n63 n137 VDD VSS XOR2_X1 
XU71 B[21] A[21] n56 VDD VSS NOR2_X1 
XU70 B[21] A[21] n58 VDD VSS NAND2_X1 
XU69 n10 n58 n59 VDD VSS NAND2_X1 
XU68 n61 n11 n60 n57 VDD VSS AOI21_X1 
XU67 n59 n57 n138 VDD VSS XOR2_X1 
XU66 n58 n56 n57 n52 VDD VSS OAI21_X1 
XU65 B[22] A[22] n53 VDD VSS AND2_X1 
XU64 B[22] A[22] n54 VDD VSS NOR2_X1 
XU63 n53 n54 n55 VDD VSS NOR2_X1 
XU62 n52 n55 n139 VDD VSS XOR2_X1 
XU61 B[23] A[23] n48 VDD VSS NOR2_X1 
XU60 B[23] A[23] n50 VDD VSS NAND2_X1 
XU59 n8 n50 n51 VDD VSS NAND2_X1 
XU58 n53 n9 n52 n49 VDD VSS AOI21_X1 
XU57 n51 n49 n140 VDD VSS XOR2_X1 
XU56 n50 n48 n49 n44 VDD VSS OAI21_X1 
XU55 B[24] A[24] n45 VDD VSS AND2_X1 
XU54 B[24] A[24] n46 VDD VSS NOR2_X1 
XU53 n45 n46 n47 VDD VSS NOR2_X1 
XU52 n44 n47 n127 VDD VSS XOR2_X1 
XU51 B[25] A[25] n40 VDD VSS NOR2_X1 
XU50 B[25] A[25] n42 VDD VSS NAND2_X1 
XU49 n6 n42 n43 VDD VSS NAND2_X1 
XU48 n45 n7 n44 n41 VDD VSS AOI21_X1 
XU47 n43 n41 n128 VDD VSS XOR2_X1 
XU46 n42 n40 n41 n36 VDD VSS OAI21_X1 
XU45 B[26] A[26] n37 VDD VSS AND2_X1 
XU1 n92 SUM[28] VDD VSS BUF_X1 
XU103 n110 SUM[22] VDD VSS BUF_X1 
XU104 n123 SUM[18] VDD VSS BUF_X1 
XU105 n133 n87 VDD VSS INV_X1 
XU106 n87 SUM[30] VDD VSS INV_X32 
XU107 n91 n89 VDD VSS INV_X1 
XU108 n89 SUM[29] VDD VSS INV_X8 
XU109 n132 n91 VDD VSS BUF_X32 
XU110 n93 n92 VDD VSS CLKBUF_X1 
XU111 n131 n93 VDD VSS BUF_X32 
XU112 n96 n94 VDD VSS INV_X1 
XU113 n94 SUM[27] VDD VSS INV_X32 
XU114 n130 n96 VDD VSS BUF_X32 
XU115 n99 n97 VDD VSS INV_X1 
XU116 n97 SUM[26] VDD VSS INV_X8 
XU117 n129 n99 VDD VSS BUF_X32 
XU118 n102 n100 VDD VSS INV_X1 
XU119 n100 SUM[25] VDD VSS INV_X8 
XU120 n128 n102 VDD VSS BUF_X32 
XU121 n105 n103 VDD VSS INV_X1 
XU122 n103 SUM[24] VDD VSS INV_X8 
XU123 n127 n105 VDD VSS BUF_X32 
XU124 n108 n106 VDD VSS INV_X1 
XU125 n106 SUM[23] VDD VSS INV_X8 
XU126 n140 n108 VDD VSS BUF_X32 
XU127 n111 n109 VDD VSS INV_X1 
XU128 n109 n110 VDD VSS INV_X4 
XU129 n139 n111 VDD VSS BUF_X32 
XU130 n114 n112 VDD VSS INV_X1 
XU131 n112 SUM[21] VDD VSS INV_X8 
XU132 n138 n114 VDD VSS BUF_X32 
XU133 n117 n115 VDD VSS INV_X1 
XU134 n115 n142 VDD VSS INV_X8 
XU135 n137 n117 VDD VSS BUF_X32 
XU136 n119 n118 VDD VSS CLKBUF_X1 
XU137 n136 n119 VDD VSS INV_X1 
XU138 n118 SUM[19] VDD VSS INV_X32 
XU139 n122 n121 VDD VSS CLKBUF_X1 
XU140 n135 n122 VDD VSS INV_X1 
XU141 n121 n123 VDD VSS INV_X32 
XU142 n125 n124 VDD VSS BUF_X1 
XU143 n134 n125 VDD VSS INV_X16 
XU144 n124 SUM[17] VDD VSS INV_X32 
XU145 n142 SUM[20] VDD VSS BUF_X1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW01_add_0 SUM[37] SUM[36] SUM[35] SUM[34] SUM[33] 
+ SUM[32] SUM[31] SUM[30] SUM[29] SUM[28] SUM[27] SUM[26] SUM[25] SUM[24] SUM[23] 
+ SUM[22] SUM[21] SUM[20] SUM[19] SUM[18] SUM[17] SUM[16] SUM[15] SUM[14] SUM[13] 
+ SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] 
+ SUM[1] SUM[0] CI CO VDD VSS B[37] B[36] B[35] B[34] B[33] B[32] B[31] B[30] B[29] 
+ B[28] B[27] B[26] B[25] B[24] B[23] B[22] B[21] B[20] B[19] B[18] B[17] B[16] 
+ B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] 
+ B[0] A[37] A[36] A[35] A[34] A[33] A[32] A[31] A[30] A[29] A[28] A[27] A[26] A[25] 
+ A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] A[13] A[12] 
+ A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU1_13 A[13] B[13] carry[13] carry[14] SUM[13] VDD VSS FA_X1 
XU1_14 A[14] B[14] carry[14] carry[15] SUM[14] VDD VSS FA_X1 
XU1_15 A[15] B[15] carry[15] carry[16] SUM[15] VDD VSS FA_X1 
XU1_16 A[16] B[16] carry[16] carry[17] SUM[16] VDD VSS FA_X1 
XU1_17 A[17] B[17] carry[17] carry[18] SUM[17] VDD VSS FA_X1 
XU1_18 A[18] B[18] carry[18] carry[19] SUM[18] VDD VSS FA_X1 
XU1_19 A[19] B[19] carry[19] carry[20] SUM[19] VDD VSS FA_X1 
XU1_20 A[20] B[20] carry[20] carry[21] n75 VDD VSS FA_X1 
XU1_21 A[21] B[21] carry[21] carry[22] n76 VDD VSS FA_X1 
XU1_22 A[22] B[22] carry[22] carry[23] n77 VDD VSS FA_X1 
XU1_23 A[23] B[23] carry[23] carry[24] n78 VDD VSS FA_X1 
XU1_24 A[24] B[24] carry[24] carry[25] n79 VDD VSS FA_X1 
XU1_25 A[25] B[25] carry[25] carry[26] n80 VDD VSS FA_X1 
XU1_26 A[26] B[26] carry[26] carry[27] n81 VDD VSS FA_X1 
XU1_27 A[27] B[27] carry[27] carry[28] n82 VDD VSS FA_X1 
XU1_28 A[28] B[28] carry[28] carry[29] n67 VDD VSS FA_X1 
XU1_29 A[29] B[29] carry[29] carry[30] n68 VDD VSS FA_X1 
XU1_30 A[30] B[30] carry[30] carry[31] n69 VDD VSS FA_X1 
XU1_31 A[31] B[31] carry[31] carry[32] n70 VDD VSS FA_X1 
XU1_32 A[32] B[32] carry[32] carry[33] n71 VDD VSS FA_X1 
XU1_33 A[33] B[33] carry[33] carry[34] n72 VDD VSS FA_X1 
XU1_34 A[34] B[34] carry[34] carry[35] n73 VDD VSS FA_X1 
XU1_35 A[35] B[35] carry[35] carry[36] n74 VDD VSS FA_X1 
XU1_36 A[36] B[36] carry[36] carry[37] n65 VDD VSS FA_X1 
XU1_37 A[37] B[37] carry[37] SYNOPSYS_UNCONNECTED_95 n66 VDD VSS FA_X1 
XU2 B[0] A[0] SUM[0] VDD VSS XOR2_X1 
XU1 B[0] A[0] n1 VDD VSS AND2_X1 
XU1_1 A[1] B[1] n1 carry[2] SUM[1] VDD VSS FA_X1 
XU1_2 A[2] B[2] carry[2] carry[3] SUM[2] VDD VSS FA_X1 
XU1_3 A[3] B[3] carry[3] carry[4] SUM[3] VDD VSS FA_X1 
XU1_4 A[4] B[4] carry[4] carry[5] SUM[4] VDD VSS FA_X1 
XU1_5 A[5] B[5] carry[5] carry[6] SUM[5] VDD VSS FA_X1 
XU1_6 A[6] B[6] carry[6] carry[7] SUM[6] VDD VSS FA_X1 
XU1_7 A[7] B[7] carry[7] carry[8] SUM[7] VDD VSS FA_X1 
XU1_8 A[8] B[8] carry[8] carry[9] SUM[8] VDD VSS FA_X1 
XU1_9 A[9] B[9] carry[9] carry[10] SUM[9] VDD VSS FA_X1 
XU1_10 A[10] B[10] carry[10] carry[11] SUM[10] VDD VSS FA_X1 
XU1_11 A[11] B[11] carry[11] carry[12] SUM[11] VDD VSS FA_X1 
XU1_12 A[12] B[12] carry[12] carry[13] SUM[12] VDD VSS FA_X1 
XU3 n3 n2 VDD VSS CLKBUF_X1 
XU4 n66 n3 VDD VSS INV_X32 
XU5 n2 SUM[37] VDD VSS INV_X32 
XU6 n6 n5 VDD VSS CLKBUF_X1 
XU7 n65 n6 VDD VSS INV_X32 
XU8 n5 SUM[36] VDD VSS INV_X32 
XU9 n11 SUM[35] VDD VSS BUF_X1 
XU10 n10 n9 VDD VSS CLKBUF_X1 
XU11 n74 n10 VDD VSS INV_X32 
XU12 n9 n11 VDD VSS INV_X32 
XU13 n13 n12 VDD VSS CLKBUF_X1 
XU14 n73 n13 VDD VSS INV_X32 
XU15 n12 SUM[34] VDD VSS INV_X32 
XU16 n18 SUM[33] VDD VSS BUF_X1 
XU17 n17 n16 VDD VSS CLKBUF_X1 
XU18 n72 n17 VDD VSS INV_X32 
XU19 n16 n18 VDD VSS INV_X32 
XU20 n22 SUM[32] VDD VSS BUF_X1 
XU21 n21 n20 VDD VSS CLKBUF_X1 
XU22 n71 n21 VDD VSS INV_X32 
XU23 n20 n22 VDD VSS INV_X32 
XU24 n26 SUM[31] VDD VSS BUF_X1 
XU25 n25 n24 VDD VSS CLKBUF_X1 
XU26 n70 n25 VDD VSS INV_X32 
XU27 n24 n26 VDD VSS INV_X32 
XU28 n28 n27 VDD VSS CLKBUF_X1 
XU29 n69 n28 VDD VSS INV_X32 
XU30 n27 SUM[30] VDD VSS INV_X32 
XU31 n31 n30 VDD VSS CLKBUF_X1 
XU32 n68 n31 VDD VSS INV_X32 
XU33 n30 SUM[29] VDD VSS INV_X32 
XU34 n34 n33 VDD VSS CLKBUF_X1 
XU35 n67 n34 VDD VSS INV_X32 
XU36 n33 SUM[28] VDD VSS INV_X32 
XU37 n37 n36 VDD VSS CLKBUF_X1 
XU38 n82 n37 VDD VSS INV_X32 
XU39 n36 SUM[27] VDD VSS INV_X32 
XU40 n40 n39 VDD VSS CLKBUF_X1 
XU41 n81 n40 VDD VSS INV_X32 
XU42 n39 SUM[26] VDD VSS INV_X32 
XU43 n43 n42 VDD VSS CLKBUF_X1 
XU44 n80 n43 VDD VSS INV_X32 
XU45 n42 SUM[25] VDD VSS INV_X32 
XU46 n48 SUM[24] VDD VSS BUF_X1 
XU47 n47 n46 VDD VSS CLKBUF_X1 
XU48 n79 n47 VDD VSS INV_X32 
XU49 n46 n48 VDD VSS INV_X32 
XU50 n52 SUM[23] VDD VSS BUF_X1 
XU51 n51 n50 VDD VSS CLKBUF_X1 
XU52 n78 n51 VDD VSS INV_X32 
XU53 n50 n52 VDD VSS INV_X32 
XU54 n56 SUM[22] VDD VSS BUF_X1 
XU55 n55 n54 VDD VSS CLKBUF_X1 
XU56 n77 n55 VDD VSS INV_X32 
XU57 n54 n56 VDD VSS INV_X32 
XU58 n60 SUM[21] VDD VSS BUF_X1 
XU59 n59 n58 VDD VSS CLKBUF_X1 
XU60 n76 n59 VDD VSS INV_X32 
XU61 n58 n60 VDD VSS INV_X32 
XU62 n64 SUM[20] VDD VSS BUF_X1 
XU63 n63 n62 VDD VSS CLKBUF_X1 
XU64 n75 n63 VDD VSS INV_X32 
XU65 n62 n64 VDD VSS INV_X32 
.ENDS

.SUBCKT gng_interp_DW01_inc_0 SUM[15] SUM[14] SUM[13] SUM[12] SUM[11] SUM[10] SUM[9] 
+ SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] A[15] A[14] A[13] 
+ A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] VDD VSS 
XU1_1_7 A[7] carry[7] carry[8] SUM[7] VDD VSS HA_X1 
XU1_1_6 A[6] carry[6] carry[7] SUM[6] VDD VSS HA_X1 
XU1_1_5 A[5] carry[5] carry[6] SUM[5] VDD VSS HA_X1 
XU1_1_4 A[4] carry[4] carry[5] SUM[4] VDD VSS HA_X1 
XU1_1_3 A[3] carry[3] carry[4] SUM[3] VDD VSS HA_X1 
XU1_1_2 A[2] carry[2] carry[3] SUM[2] VDD VSS HA_X1 
XU1_1_1 A[1] A[0] carry[2] SUM[1] VDD VSS HA_X1 
XU1 carry[15] SUM[15] VDD VSS INV_X1 
XU1_1_14 A[14] carry[14] carry[15] SUM[14] VDD VSS HA_X1 
XU1_1_13 A[13] carry[13] carry[14] SUM[13] VDD VSS HA_X1 
XU1_1_12 A[12] carry[12] carry[13] SUM[12] VDD VSS HA_X1 
XU1_1_11 A[11] carry[11] carry[12] SUM[11] VDD VSS HA_X1 
XU1_1_10 A[10] carry[10] carry[11] SUM[10] VDD VSS HA_X1 
XU1_1_9 A[9] carry[9] carry[10] SUM[9] VDD VSS HA_X1 
XU1_1_8 A[8] carry[8] carry[9] SUM[8] VDD VSS HA_X1 
.ENDS

.SUBCKT gng_interp_DW01_add_1 SUM[17] SUM[16] SUM[15] SUM[14] SUM[13] SUM[12] SUM[11] 
+ SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
+ CI CO B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] 
+ B[4] B[3] B[2] B[1] B[0] A[17] A[16] A[15] A[14] A[13] A[12] A[11] A[10] A[9] 
+ A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] VDD VSS 
XU4 A[0] B[0] A[1] B[1] n3 VDD VSS OAI211_X1 
XU3 n3 n2 n1 carry[2] VDD VSS OAI21_X1 
XU2 B[1] n1 VDD VSS INV_X1 
XU1 A[1] n2 VDD VSS INV_X1 
XU1_2 A[2] B[2] carry[2] carry[3] n74 VDD VSS FA_X1 
XU1_3 A[3] B[3] carry[3] carry[4] n75 VDD VSS FA_X1 
XU1_4 A[4] B[4] carry[4] carry[5] n66 VDD VSS FA_X1 
XU1_5 A[5] B[5] carry[5] carry[6] n67 VDD VSS FA_X1 
XU1_6 A[6] B[6] carry[6] carry[7] n68 VDD VSS FA_X1 
XU1_7 A[7] B[7] carry[7] carry[8] n69 VDD VSS FA_X1 
XU1_8 A[8] B[8] carry[8] carry[9] n70 VDD VSS FA_X1 
XU1_9 A[9] B[9] carry[9] carry[10] n71 VDD VSS FA_X1 
XU1_10 A[10] B[10] carry[10] carry[11] n72 VDD VSS FA_X1 
XU1_11 A[11] B[11] carry[11] carry[12] n73 VDD VSS FA_X1 
XU1_12 A[12] B[12] carry[12] carry[13] n60 VDD VSS FA_X1 
XU1_13 A[13] B[13] carry[13] carry[14] n61 VDD VSS FA_X1 
XU1_14 A[14] B[14] carry[14] carry[15] n62 VDD VSS FA_X1 
XU1_15 A[15] B[15] carry[15] carry[16] n63 VDD VSS FA_X1 
XU1_16 A[16] B[16] carry[16] carry[17] n64 VDD VSS FA_X1 
XU1_17 A[17] B[17] carry[17] SYNOPSYS_UNCONNECTED_44 n65 VDD VSS FA_X1 
XU5 n7 SUM[17] VDD VSS BUF_X1 
XU6 n6 n5 VDD VSS CLKBUF_X1 
XU7 n65 n6 VDD VSS INV_X32 
XU8 n5 n7 VDD VSS INV_X32 
XU9 n11 SUM[16] VDD VSS BUF_X1 
XU10 n10 n9 VDD VSS CLKBUF_X1 
XU11 n64 n10 VDD VSS INV_X32 
XU12 n9 n11 VDD VSS INV_X32 
XU13 n15 SUM[15] VDD VSS BUF_X1 
XU14 n14 n13 VDD VSS CLKBUF_X1 
XU15 n63 n14 VDD VSS INV_X32 
XU16 n13 n15 VDD VSS INV_X32 
XU17 n62 n16 VDD VSS CLKBUF_X1 
XU18 n18 n17 VDD VSS CLKBUF_X1 
XU19 n16 n18 VDD VSS INV_X32 
XU20 n17 SUM[14] VDD VSS INV_X32 
XU21 n23 SUM[13] VDD VSS CLKBUF_X1 
XU22 n22 n21 VDD VSS CLKBUF_X1 
XU23 n61 n22 VDD VSS INV_X32 
XU24 n21 n23 VDD VSS INV_X32 
XU25 n27 SUM[12] VDD VSS BUF_X1 
XU26 n26 n25 VDD VSS CLKBUF_X1 
XU27 n60 n26 VDD VSS INV_X32 
XU28 n25 n27 VDD VSS INV_X32 
XU29 n73 n28 VDD VSS CLKBUF_X1 
XU30 n30 n29 VDD VSS CLKBUF_X1 
XU31 n28 n30 VDD VSS INV_X32 
XU32 n29 SUM[11] VDD VSS INV_X32 
XU33 n33 n32 VDD VSS CLKBUF_X1 
XU34 n72 n33 VDD VSS INV_X32 
XU35 n32 SUM[10] VDD VSS INV_X32 
XU36 n36 n35 VDD VSS BUF_X1 
XU37 n71 n36 VDD VSS INV_X32 
XU38 n35 SUM[9] VDD VSS INV_X32 
XU39 n39 n38 VDD VSS BUF_X1 
XU40 n70 n39 VDD VSS INV_X32 
XU41 n38 SUM[8] VDD VSS INV_X32 
XU42 n42 n41 VDD VSS CLKBUF_X1 
XU43 n69 n42 VDD VSS INV_X32 
XU44 n41 SUM[7] VDD VSS INV_X16 
XU45 n47 SUM[6] VDD VSS BUF_X1 
XU46 n46 n45 VDD VSS CLKBUF_X1 
XU47 n68 n46 VDD VSS INV_X32 
XU48 n45 n47 VDD VSS INV_X32 
XU49 n49 n48 VDD VSS CLKBUF_X1 
XU50 n67 n49 VDD VSS INV_X32 
XU51 n48 SUM[5] VDD VSS INV_X32 
XU52 n52 n51 VDD VSS CLKBUF_X1 
XU53 n66 n52 VDD VSS INV_X32 
XU54 n51 SUM[4] VDD VSS INV_X32 
XU55 n55 n54 VDD VSS BUF_X1 
XU56 n75 n55 VDD VSS INV_X32 
XU57 n54 SUM[3] VDD VSS INV_X32 
XU58 n58 n57 VDD VSS BUF_X1 
XU59 n74 n58 VDD VSS INV_X32 
XU60 n57 SUM[2] VDD VSS INV_X32 
.ENDS

.SUBCKT gng_smul_16_18_DW02_mult_0 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] 
+ PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] PRODUCT[1] 
+ PRODUCT[0] TC VDD VSS B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] 
+ B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] 
+ A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XS2_14_3 ab_14__3_ CARRYB_13__3_ SUMB_13__4_ CARRYB_14__3_ SUMB_14__3_ VDD VSS FA_X1 
XS2_14_2 ab_14__2_ CARRYB_13__2_ SUMB_13__3_ CARRYB_14__2_ SUMB_14__2_ VDD VSS FA_X1 
XS2_14_1 ab_14__1_ CARRYB_13__1_ SUMB_13__2_ CARRYB_14__1_ SUMB_14__1_ VDD VSS FA_X1 
XS1_14_0 ab_14__0_ CARRYB_13__0_ SUMB_13__1_ CARRYB_14__0_ PRODUCT[14] VDD VSS FA_X1 
XS14_17 n1 n85 ab_15__17_ CARRYB_15__17_ SUMB_15__17_ VDD VSS FA_X1 
XS5_16 ab_15__16_ CARRYB_14__16_ ab_14__17_ CARRYB_15__16_ SUMB_15__16_ VDD VSS FA_X1 
XS4_15 ab_15__15_ CARRYB_14__15_ SUMB_14__16_ CARRYB_15__15_ SUMB_15__15_ VDD VSS FA_X1 
XS4_14 ab_15__14_ CARRYB_14__14_ SUMB_14__15_ CARRYB_15__14_ SUMB_15__14_ VDD VSS FA_X1 
XS4_13 ab_15__13_ CARRYB_14__13_ SUMB_14__14_ CARRYB_15__13_ SUMB_15__13_ VDD VSS FA_X1 
XS4_12 ab_15__12_ CARRYB_14__12_ SUMB_14__13_ CARRYB_15__12_ SUMB_15__12_ VDD VSS FA_X1 
XS4_11 ab_15__11_ CARRYB_14__11_ SUMB_14__12_ CARRYB_15__11_ SUMB_15__11_ VDD VSS FA_X1 
XS4_10 ab_15__10_ CARRYB_14__10_ SUMB_14__11_ CARRYB_15__10_ SUMB_15__10_ VDD VSS FA_X1 
XS4_9 ab_15__9_ CARRYB_14__9_ SUMB_14__10_ CARRYB_15__9_ SUMB_15__9_ VDD VSS FA_X1 
XS4_8 ab_15__8_ CARRYB_14__8_ SUMB_14__9_ CARRYB_15__8_ SUMB_15__8_ VDD VSS FA_X1 
XS4_7 ab_15__7_ CARRYB_14__7_ SUMB_14__8_ CARRYB_15__7_ SUMB_15__7_ VDD VSS FA_X1 
XS4_6 ab_15__6_ CARRYB_14__6_ SUMB_14__7_ CARRYB_15__6_ SUMB_15__6_ VDD VSS FA_X1 
XS4_5 ab_15__5_ CARRYB_14__5_ SUMB_14__6_ CARRYB_15__5_ SUMB_15__5_ VDD VSS FA_X1 
XS4_4 ab_15__4_ CARRYB_14__4_ SUMB_14__5_ CARRYB_15__4_ SUMB_15__4_ VDD VSS FA_X1 
XS4_3 ab_15__3_ CARRYB_14__3_ SUMB_14__4_ CARRYB_15__3_ SUMB_15__3_ VDD VSS FA_X1 
XS4_2 ab_15__2_ CARRYB_14__2_ SUMB_14__3_ CARRYB_15__2_ SUMB_15__2_ VDD VSS FA_X1 
XS4_1 ab_15__1_ CARRYB_14__1_ SUMB_14__2_ CARRYB_15__1_ SUMB_15__1_ VDD VSS FA_X1 
XS4_0 ab_15__0_ CARRYB_14__0_ SUMB_14__1_ CARRYB_15__0_ SUMB_15__0_ VDD VSS FA_X1 
XS14_17_0 B[17] CARRYB_15__1_ SUMB_15__2_ A2_16_ A1_15_ VDD VSS FA_X1 
XS2_9_11 ab_9__11_ CARRYB_8__11_ SUMB_8__12_ CARRYB_9__11_ SUMB_9__11_ VDD VSS FA_X1 
XS2_9_10 ab_9__10_ CARRYB_8__10_ SUMB_8__11_ CARRYB_9__10_ SUMB_9__10_ VDD VSS FA_X1 
XS2_9_9 ab_9__9_ CARRYB_8__9_ SUMB_8__10_ CARRYB_9__9_ SUMB_9__9_ VDD VSS FA_X1 
XS2_9_8 ab_9__8_ CARRYB_8__8_ SUMB_8__9_ CARRYB_9__8_ SUMB_9__8_ VDD VSS FA_X1 
XS2_9_7 ab_9__7_ CARRYB_8__7_ SUMB_8__8_ CARRYB_9__7_ SUMB_9__7_ VDD VSS FA_X1 
XS2_9_6 ab_9__6_ CARRYB_8__6_ SUMB_8__7_ CARRYB_9__6_ SUMB_9__6_ VDD VSS FA_X1 
XS2_9_5 ab_9__5_ CARRYB_8__5_ SUMB_8__6_ CARRYB_9__5_ SUMB_9__5_ VDD VSS FA_X1 
XS2_9_4 ab_9__4_ CARRYB_8__4_ SUMB_8__5_ CARRYB_9__4_ SUMB_9__4_ VDD VSS FA_X1 
XS2_9_3 ab_9__3_ CARRYB_8__3_ SUMB_8__4_ CARRYB_9__3_ SUMB_9__3_ VDD VSS FA_X1 
XS2_9_2 ab_9__2_ CARRYB_8__2_ SUMB_8__3_ CARRYB_9__2_ SUMB_9__2_ VDD VSS FA_X1 
XS2_9_1 ab_9__1_ CARRYB_8__1_ SUMB_8__2_ CARRYB_9__1_ SUMB_9__1_ VDD VSS FA_X1 
XS1_9_0 ab_9__0_ CARRYB_8__0_ SUMB_8__1_ CARRYB_9__0_ PRODUCT[9] VDD VSS FA_X1 
XS3_10_16 ab_10__16_ CARRYB_9__16_ ab_9__17_ CARRYB_10__16_ SUMB_10__16_ VDD VSS FA_X1 
XS2_10_15 ab_10__15_ CARRYB_9__15_ SUMB_9__16_ CARRYB_10__15_ SUMB_10__15_ VDD VSS FA_X1 
XS2_10_14 ab_10__14_ CARRYB_9__14_ SUMB_9__15_ CARRYB_10__14_ SUMB_10__14_ VDD VSS FA_X1 
XS2_10_13 ab_10__13_ CARRYB_9__13_ SUMB_9__14_ CARRYB_10__13_ SUMB_10__13_ VDD VSS FA_X1 
XS2_10_12 ab_10__12_ CARRYB_9__12_ SUMB_9__13_ CARRYB_10__12_ SUMB_10__12_ VDD VSS FA_X1 
XS2_10_11 ab_10__11_ CARRYB_9__11_ SUMB_9__12_ CARRYB_10__11_ SUMB_10__11_ VDD VSS FA_X1 
XS2_10_10 ab_10__10_ CARRYB_9__10_ SUMB_9__11_ CARRYB_10__10_ SUMB_10__10_ VDD VSS FA_X1 
XS2_10_9 ab_10__9_ CARRYB_9__9_ SUMB_9__10_ CARRYB_10__9_ SUMB_10__9_ VDD VSS FA_X1 
XS2_10_8 ab_10__8_ CARRYB_9__8_ SUMB_9__9_ CARRYB_10__8_ SUMB_10__8_ VDD VSS FA_X1 
XS2_10_7 ab_10__7_ CARRYB_9__7_ SUMB_9__8_ CARRYB_10__7_ SUMB_10__7_ VDD VSS FA_X1 
XS2_10_6 ab_10__6_ CARRYB_9__6_ SUMB_9__7_ CARRYB_10__6_ SUMB_10__6_ VDD VSS FA_X1 
XS2_10_5 ab_10__5_ CARRYB_9__5_ SUMB_9__6_ CARRYB_10__5_ SUMB_10__5_ VDD VSS FA_X1 
XS2_10_4 ab_10__4_ CARRYB_9__4_ SUMB_9__5_ CARRYB_10__4_ SUMB_10__4_ VDD VSS FA_X1 
XS2_10_3 ab_10__3_ CARRYB_9__3_ SUMB_9__4_ CARRYB_10__3_ SUMB_10__3_ VDD VSS FA_X1 
XS2_10_2 ab_10__2_ CARRYB_9__2_ SUMB_9__3_ CARRYB_10__2_ SUMB_10__2_ VDD VSS FA_X1 
XS2_10_1 ab_10__1_ CARRYB_9__1_ SUMB_9__2_ CARRYB_10__1_ SUMB_10__1_ VDD VSS FA_X1 
XS1_10_0 ab_10__0_ CARRYB_9__0_ SUMB_9__1_ CARRYB_10__0_ PRODUCT[10] VDD VSS FA_X1 
XS3_11_16 ab_11__16_ CARRYB_10__16_ ab_10__17_ CARRYB_11__16_ SUMB_11__16_ VDD VSS FA_X1 
XS2_11_15 ab_11__15_ CARRYB_10__15_ SUMB_10__16_ CARRYB_11__15_ SUMB_11__15_ VDD 
+ VSS FA_X1 
XS2_11_14 ab_11__14_ CARRYB_10__14_ SUMB_10__15_ CARRYB_11__14_ SUMB_11__14_ VDD 
+ VSS FA_X1 
XS2_11_13 ab_11__13_ CARRYB_10__13_ SUMB_10__14_ CARRYB_11__13_ SUMB_11__13_ VDD 
+ VSS FA_X1 
XS2_11_12 ab_11__12_ CARRYB_10__12_ SUMB_10__13_ CARRYB_11__12_ SUMB_11__12_ VDD 
+ VSS FA_X1 
XS2_11_11 ab_11__11_ CARRYB_10__11_ SUMB_10__12_ CARRYB_11__11_ SUMB_11__11_ VDD 
+ VSS FA_X1 
XS2_11_10 ab_11__10_ CARRYB_10__10_ SUMB_10__11_ CARRYB_11__10_ SUMB_11__10_ VDD 
+ VSS FA_X1 
XS2_11_9 ab_11__9_ CARRYB_10__9_ SUMB_10__10_ CARRYB_11__9_ SUMB_11__9_ VDD VSS FA_X1 
XS2_11_8 ab_11__8_ CARRYB_10__8_ SUMB_10__9_ CARRYB_11__8_ SUMB_11__8_ VDD VSS FA_X1 
XS2_11_7 ab_11__7_ CARRYB_10__7_ SUMB_10__8_ CARRYB_11__7_ SUMB_11__7_ VDD VSS FA_X1 
XS2_11_6 ab_11__6_ CARRYB_10__6_ SUMB_10__7_ CARRYB_11__6_ SUMB_11__6_ VDD VSS FA_X1 
XS2_11_5 ab_11__5_ CARRYB_10__5_ SUMB_10__6_ CARRYB_11__5_ SUMB_11__5_ VDD VSS FA_X1 
XS2_11_4 ab_11__4_ CARRYB_10__4_ SUMB_10__5_ CARRYB_11__4_ SUMB_11__4_ VDD VSS FA_X1 
XS2_11_3 ab_11__3_ CARRYB_10__3_ SUMB_10__4_ CARRYB_11__3_ SUMB_11__3_ VDD VSS FA_X1 
XS2_11_2 ab_11__2_ CARRYB_10__2_ SUMB_10__3_ CARRYB_11__2_ SUMB_11__2_ VDD VSS FA_X1 
XS2_11_1 ab_11__1_ CARRYB_10__1_ SUMB_10__2_ CARRYB_11__1_ SUMB_11__1_ VDD VSS FA_X1 
XS1_11_0 ab_11__0_ CARRYB_10__0_ SUMB_10__1_ CARRYB_11__0_ PRODUCT[11] VDD VSS FA_X1 
XS3_12_16 ab_12__16_ CARRYB_11__16_ ab_11__17_ CARRYB_12__16_ SUMB_12__16_ VDD VSS FA_X1 
XS2_12_15 ab_12__15_ CARRYB_11__15_ SUMB_11__16_ CARRYB_12__15_ SUMB_12__15_ VDD 
+ VSS FA_X1 
XS2_12_14 ab_12__14_ CARRYB_11__14_ SUMB_11__15_ CARRYB_12__14_ SUMB_12__14_ VDD 
+ VSS FA_X1 
XS2_12_13 ab_12__13_ CARRYB_11__13_ SUMB_11__14_ CARRYB_12__13_ SUMB_12__13_ VDD 
+ VSS FA_X1 
XS2_12_12 ab_12__12_ CARRYB_11__12_ SUMB_11__13_ CARRYB_12__12_ SUMB_12__12_ VDD 
+ VSS FA_X1 
XS2_12_11 ab_12__11_ CARRYB_11__11_ SUMB_11__12_ CARRYB_12__11_ SUMB_12__11_ VDD 
+ VSS FA_X1 
XS2_12_10 ab_12__10_ CARRYB_11__10_ SUMB_11__11_ CARRYB_12__10_ SUMB_12__10_ VDD 
+ VSS FA_X1 
XS2_12_9 ab_12__9_ CARRYB_11__9_ SUMB_11__10_ CARRYB_12__9_ SUMB_12__9_ VDD VSS FA_X1 
XS2_12_8 ab_12__8_ CARRYB_11__8_ SUMB_11__9_ CARRYB_12__8_ SUMB_12__8_ VDD VSS FA_X1 
XS2_12_7 ab_12__7_ CARRYB_11__7_ SUMB_11__8_ CARRYB_12__7_ SUMB_12__7_ VDD VSS FA_X1 
XS2_12_6 ab_12__6_ CARRYB_11__6_ SUMB_11__7_ CARRYB_12__6_ SUMB_12__6_ VDD VSS FA_X1 
XS2_12_5 ab_12__5_ CARRYB_11__5_ SUMB_11__6_ CARRYB_12__5_ SUMB_12__5_ VDD VSS FA_X1 
XS2_12_4 ab_12__4_ CARRYB_11__4_ SUMB_11__5_ CARRYB_12__4_ SUMB_12__4_ VDD VSS FA_X1 
XS2_12_3 ab_12__3_ CARRYB_11__3_ SUMB_11__4_ CARRYB_12__3_ SUMB_12__3_ VDD VSS FA_X1 
XS2_12_2 ab_12__2_ CARRYB_11__2_ SUMB_11__3_ CARRYB_12__2_ SUMB_12__2_ VDD VSS FA_X1 
XS2_12_1 ab_12__1_ CARRYB_11__1_ SUMB_11__2_ CARRYB_12__1_ SUMB_12__1_ VDD VSS FA_X1 
XS1_12_0 ab_12__0_ CARRYB_11__0_ SUMB_11__1_ CARRYB_12__0_ PRODUCT[12] VDD VSS FA_X1 
XS3_13_16 ab_13__16_ CARRYB_12__16_ ab_12__17_ CARRYB_13__16_ SUMB_13__16_ VDD VSS FA_X1 
XS2_13_15 ab_13__15_ CARRYB_12__15_ SUMB_12__16_ CARRYB_13__15_ SUMB_13__15_ VDD 
+ VSS FA_X1 
XS2_13_14 ab_13__14_ CARRYB_12__14_ SUMB_12__15_ CARRYB_13__14_ SUMB_13__14_ VDD 
+ VSS FA_X1 
XS2_13_13 ab_13__13_ CARRYB_12__13_ SUMB_12__14_ CARRYB_13__13_ SUMB_13__13_ VDD 
+ VSS FA_X1 
XS2_13_12 ab_13__12_ CARRYB_12__12_ SUMB_12__13_ CARRYB_13__12_ SUMB_13__12_ VDD 
+ VSS FA_X1 
XS2_13_11 ab_13__11_ CARRYB_12__11_ SUMB_12__12_ CARRYB_13__11_ SUMB_13__11_ VDD 
+ VSS FA_X1 
XS2_13_10 ab_13__10_ CARRYB_12__10_ SUMB_12__11_ CARRYB_13__10_ SUMB_13__10_ VDD 
+ VSS FA_X1 
XS2_13_9 ab_13__9_ CARRYB_12__9_ SUMB_12__10_ CARRYB_13__9_ SUMB_13__9_ VDD VSS FA_X1 
XS2_13_8 ab_13__8_ CARRYB_12__8_ SUMB_12__9_ CARRYB_13__8_ SUMB_13__8_ VDD VSS FA_X1 
XS2_13_7 ab_13__7_ CARRYB_12__7_ SUMB_12__8_ CARRYB_13__7_ SUMB_13__7_ VDD VSS FA_X1 
XS2_13_6 ab_13__6_ CARRYB_12__6_ SUMB_12__7_ CARRYB_13__6_ SUMB_13__6_ VDD VSS FA_X1 
XS2_13_5 ab_13__5_ CARRYB_12__5_ SUMB_12__6_ CARRYB_13__5_ SUMB_13__5_ VDD VSS FA_X1 
XS2_13_4 ab_13__4_ CARRYB_12__4_ SUMB_12__5_ CARRYB_13__4_ SUMB_13__4_ VDD VSS FA_X1 
XS2_13_3 ab_13__3_ CARRYB_12__3_ SUMB_12__4_ CARRYB_13__3_ SUMB_13__3_ VDD VSS FA_X1 
XS2_13_2 ab_13__2_ CARRYB_12__2_ SUMB_12__3_ CARRYB_13__2_ SUMB_13__2_ VDD VSS FA_X1 
XS2_13_1 ab_13__1_ CARRYB_12__1_ SUMB_12__2_ CARRYB_13__1_ SUMB_13__1_ VDD VSS FA_X1 
XS1_13_0 ab_13__0_ CARRYB_12__0_ SUMB_12__1_ CARRYB_13__0_ PRODUCT[13] VDD VSS FA_X1 
XS3_14_16 ab_14__16_ CARRYB_13__16_ ab_13__17_ CARRYB_14__16_ SUMB_14__16_ VDD VSS FA_X1 
XS2_14_15 ab_14__15_ CARRYB_13__15_ SUMB_13__16_ CARRYB_14__15_ SUMB_14__15_ VDD 
+ VSS FA_X1 
XS2_14_14 ab_14__14_ CARRYB_13__14_ SUMB_13__15_ CARRYB_14__14_ SUMB_14__14_ VDD 
+ VSS FA_X1 
XS2_14_13 ab_14__13_ CARRYB_13__13_ SUMB_13__14_ CARRYB_14__13_ SUMB_14__13_ VDD 
+ VSS FA_X1 
XS2_14_12 ab_14__12_ CARRYB_13__12_ SUMB_13__13_ CARRYB_14__12_ SUMB_14__12_ VDD 
+ VSS FA_X1 
XS2_14_11 ab_14__11_ CARRYB_13__11_ SUMB_13__12_ CARRYB_14__11_ SUMB_14__11_ VDD 
+ VSS FA_X1 
XS2_14_10 ab_14__10_ CARRYB_13__10_ SUMB_13__11_ CARRYB_14__10_ SUMB_14__10_ VDD 
+ VSS FA_X1 
XS2_14_9 ab_14__9_ CARRYB_13__9_ SUMB_13__10_ CARRYB_14__9_ SUMB_14__9_ VDD VSS FA_X1 
XS2_14_8 ab_14__8_ CARRYB_13__8_ SUMB_13__9_ CARRYB_14__8_ SUMB_14__8_ VDD VSS FA_X1 
XS2_14_7 ab_14__7_ CARRYB_13__7_ SUMB_13__8_ CARRYB_14__7_ SUMB_14__7_ VDD VSS FA_X1 
XS2_14_6 ab_14__6_ CARRYB_13__6_ SUMB_13__7_ CARRYB_14__6_ SUMB_14__6_ VDD VSS FA_X1 
XS2_14_5 ab_14__5_ CARRYB_13__5_ SUMB_13__6_ CARRYB_14__5_ SUMB_14__5_ VDD VSS FA_X1 
XS2_14_4 ab_14__4_ CARRYB_13__4_ SUMB_13__5_ CARRYB_14__4_ SUMB_14__4_ VDD VSS FA_X1 
XS2_3_2 ab_3__2_ CARRYB_2__2_ SUMB_2__3_ CARRYB_3__2_ SUMB_3__2_ VDD VSS FA_X1 
XS2_3_1 ab_3__1_ CARRYB_2__1_ SUMB_2__2_ CARRYB_3__1_ SUMB_3__1_ VDD VSS FA_X1 
XS1_3_0 ab_3__0_ CARRYB_2__0_ SUMB_2__1_ CARRYB_3__0_ PRODUCT[3] VDD VSS FA_X1 
XS3_4_16 ab_4__16_ CARRYB_3__16_ ab_3__17_ CARRYB_4__16_ SUMB_4__16_ VDD VSS FA_X1 
XS2_4_15 ab_4__15_ CARRYB_3__15_ SUMB_3__16_ CARRYB_4__15_ SUMB_4__15_ VDD VSS FA_X1 
XS2_4_14 ab_4__14_ CARRYB_3__14_ SUMB_3__15_ CARRYB_4__14_ SUMB_4__14_ VDD VSS FA_X1 
XS2_4_13 ab_4__13_ CARRYB_3__13_ SUMB_3__14_ CARRYB_4__13_ SUMB_4__13_ VDD VSS FA_X1 
XS2_4_12 ab_4__12_ CARRYB_3__12_ SUMB_3__13_ CARRYB_4__12_ SUMB_4__12_ VDD VSS FA_X1 
XS2_4_11 ab_4__11_ CARRYB_3__11_ SUMB_3__12_ CARRYB_4__11_ SUMB_4__11_ VDD VSS FA_X1 
XS2_4_10 ab_4__10_ CARRYB_3__10_ SUMB_3__11_ CARRYB_4__10_ SUMB_4__10_ VDD VSS FA_X1 
XS2_4_9 ab_4__9_ CARRYB_3__9_ SUMB_3__10_ CARRYB_4__9_ SUMB_4__9_ VDD VSS FA_X1 
XS2_4_8 ab_4__8_ CARRYB_3__8_ SUMB_3__9_ CARRYB_4__8_ SUMB_4__8_ VDD VSS FA_X1 
XS2_4_7 ab_4__7_ CARRYB_3__7_ SUMB_3__8_ CARRYB_4__7_ SUMB_4__7_ VDD VSS FA_X1 
XS2_4_6 ab_4__6_ CARRYB_3__6_ SUMB_3__7_ CARRYB_4__6_ SUMB_4__6_ VDD VSS FA_X1 
XS2_4_5 ab_4__5_ CARRYB_3__5_ SUMB_3__6_ CARRYB_4__5_ SUMB_4__5_ VDD VSS FA_X1 
XS2_4_4 ab_4__4_ CARRYB_3__4_ SUMB_3__5_ CARRYB_4__4_ SUMB_4__4_ VDD VSS FA_X1 
XS2_4_3 ab_4__3_ CARRYB_3__3_ SUMB_3__4_ CARRYB_4__3_ SUMB_4__3_ VDD VSS FA_X1 
XS2_4_2 ab_4__2_ CARRYB_3__2_ SUMB_3__3_ CARRYB_4__2_ SUMB_4__2_ VDD VSS FA_X1 
XS2_4_1 ab_4__1_ CARRYB_3__1_ SUMB_3__2_ CARRYB_4__1_ SUMB_4__1_ VDD VSS FA_X1 
XS1_4_0 ab_4__0_ CARRYB_3__0_ SUMB_3__1_ CARRYB_4__0_ PRODUCT[4] VDD VSS FA_X1 
XS3_5_16 ab_5__16_ CARRYB_4__16_ ab_4__17_ CARRYB_5__16_ SUMB_5__16_ VDD VSS FA_X1 
XS2_5_15 ab_5__15_ CARRYB_4__15_ SUMB_4__16_ CARRYB_5__15_ SUMB_5__15_ VDD VSS FA_X1 
XS2_5_14 ab_5__14_ CARRYB_4__14_ SUMB_4__15_ CARRYB_5__14_ SUMB_5__14_ VDD VSS FA_X1 
XS2_5_13 ab_5__13_ CARRYB_4__13_ SUMB_4__14_ CARRYB_5__13_ SUMB_5__13_ VDD VSS FA_X1 
XS2_5_12 ab_5__12_ CARRYB_4__12_ SUMB_4__13_ CARRYB_5__12_ SUMB_5__12_ VDD VSS FA_X1 
XS2_5_11 ab_5__11_ CARRYB_4__11_ SUMB_4__12_ CARRYB_5__11_ SUMB_5__11_ VDD VSS FA_X1 
XS2_5_10 ab_5__10_ CARRYB_4__10_ SUMB_4__11_ CARRYB_5__10_ SUMB_5__10_ VDD VSS FA_X1 
XS2_5_9 ab_5__9_ CARRYB_4__9_ SUMB_4__10_ CARRYB_5__9_ SUMB_5__9_ VDD VSS FA_X1 
XS2_5_8 ab_5__8_ CARRYB_4__8_ SUMB_4__9_ CARRYB_5__8_ SUMB_5__8_ VDD VSS FA_X1 
XS2_5_7 ab_5__7_ CARRYB_4__7_ SUMB_4__8_ CARRYB_5__7_ SUMB_5__7_ VDD VSS FA_X1 
XS2_5_6 ab_5__6_ CARRYB_4__6_ SUMB_4__7_ CARRYB_5__6_ SUMB_5__6_ VDD VSS FA_X1 
XS2_5_5 ab_5__5_ CARRYB_4__5_ SUMB_4__6_ CARRYB_5__5_ SUMB_5__5_ VDD VSS FA_X1 
XS2_5_4 ab_5__4_ CARRYB_4__4_ SUMB_4__5_ CARRYB_5__4_ SUMB_5__4_ VDD VSS FA_X1 
XS2_5_3 ab_5__3_ CARRYB_4__3_ SUMB_4__4_ CARRYB_5__3_ SUMB_5__3_ VDD VSS FA_X1 
XS2_5_2 ab_5__2_ CARRYB_4__2_ SUMB_4__3_ CARRYB_5__2_ SUMB_5__2_ VDD VSS FA_X1 
XS2_5_1 ab_5__1_ CARRYB_4__1_ SUMB_4__2_ CARRYB_5__1_ SUMB_5__1_ VDD VSS FA_X1 
XS1_5_0 ab_5__0_ CARRYB_4__0_ SUMB_4__1_ CARRYB_5__0_ PRODUCT[5] VDD VSS FA_X1 
XS3_6_16 ab_6__16_ CARRYB_5__16_ ab_5__17_ CARRYB_6__16_ SUMB_6__16_ VDD VSS FA_X1 
XS2_6_15 ab_6__15_ CARRYB_5__15_ SUMB_5__16_ CARRYB_6__15_ SUMB_6__15_ VDD VSS FA_X1 
XS2_6_14 ab_6__14_ CARRYB_5__14_ SUMB_5__15_ CARRYB_6__14_ SUMB_6__14_ VDD VSS FA_X1 
XS2_6_13 ab_6__13_ CARRYB_5__13_ SUMB_5__14_ CARRYB_6__13_ SUMB_6__13_ VDD VSS FA_X1 
XS2_6_12 ab_6__12_ CARRYB_5__12_ SUMB_5__13_ CARRYB_6__12_ SUMB_6__12_ VDD VSS FA_X1 
XS2_6_11 ab_6__11_ CARRYB_5__11_ SUMB_5__12_ CARRYB_6__11_ SUMB_6__11_ VDD VSS FA_X1 
XS2_6_10 ab_6__10_ CARRYB_5__10_ SUMB_5__11_ CARRYB_6__10_ SUMB_6__10_ VDD VSS FA_X1 
XS2_6_9 ab_6__9_ CARRYB_5__9_ SUMB_5__10_ CARRYB_6__9_ SUMB_6__9_ VDD VSS FA_X1 
XS2_6_8 ab_6__8_ CARRYB_5__8_ SUMB_5__9_ CARRYB_6__8_ SUMB_6__8_ VDD VSS FA_X1 
XS2_6_7 ab_6__7_ CARRYB_5__7_ SUMB_5__8_ CARRYB_6__7_ SUMB_6__7_ VDD VSS FA_X1 
XS2_6_6 ab_6__6_ CARRYB_5__6_ SUMB_5__7_ CARRYB_6__6_ SUMB_6__6_ VDD VSS FA_X1 
XS2_6_5 ab_6__5_ CARRYB_5__5_ SUMB_5__6_ CARRYB_6__5_ SUMB_6__5_ VDD VSS FA_X1 
XS2_6_4 ab_6__4_ CARRYB_5__4_ SUMB_5__5_ CARRYB_6__4_ SUMB_6__4_ VDD VSS FA_X1 
XS2_6_3 ab_6__3_ CARRYB_5__3_ SUMB_5__4_ CARRYB_6__3_ SUMB_6__3_ VDD VSS FA_X1 
XS2_6_2 ab_6__2_ CARRYB_5__2_ SUMB_5__3_ CARRYB_6__2_ SUMB_6__2_ VDD VSS FA_X1 
XS2_6_1 ab_6__1_ CARRYB_5__1_ SUMB_5__2_ CARRYB_6__1_ SUMB_6__1_ VDD VSS FA_X1 
XS1_6_0 ab_6__0_ CARRYB_5__0_ SUMB_5__1_ CARRYB_6__0_ PRODUCT[6] VDD VSS FA_X1 
XS3_7_16 ab_7__16_ CARRYB_6__16_ ab_6__17_ CARRYB_7__16_ SUMB_7__16_ VDD VSS FA_X1 
XS2_7_15 ab_7__15_ CARRYB_6__15_ SUMB_6__16_ CARRYB_7__15_ SUMB_7__15_ VDD VSS FA_X1 
XS2_7_14 ab_7__14_ CARRYB_6__14_ SUMB_6__15_ CARRYB_7__14_ SUMB_7__14_ VDD VSS FA_X1 
XS2_7_13 ab_7__13_ CARRYB_6__13_ SUMB_6__14_ CARRYB_7__13_ SUMB_7__13_ VDD VSS FA_X1 
XS2_7_12 ab_7__12_ CARRYB_6__12_ SUMB_6__13_ CARRYB_7__12_ SUMB_7__12_ VDD VSS FA_X1 
XS2_7_11 ab_7__11_ CARRYB_6__11_ SUMB_6__12_ CARRYB_7__11_ SUMB_7__11_ VDD VSS FA_X1 
XS2_7_10 ab_7__10_ CARRYB_6__10_ SUMB_6__11_ CARRYB_7__10_ SUMB_7__10_ VDD VSS FA_X1 
XS2_7_9 ab_7__9_ CARRYB_6__9_ SUMB_6__10_ CARRYB_7__9_ SUMB_7__9_ VDD VSS FA_X1 
XS2_7_8 ab_7__8_ CARRYB_6__8_ SUMB_6__9_ CARRYB_7__8_ SUMB_7__8_ VDD VSS FA_X1 
XS2_7_7 ab_7__7_ CARRYB_6__7_ SUMB_6__8_ CARRYB_7__7_ SUMB_7__7_ VDD VSS FA_X1 
XS2_7_6 ab_7__6_ CARRYB_6__6_ SUMB_6__7_ CARRYB_7__6_ SUMB_7__6_ VDD VSS FA_X1 
XS2_7_5 ab_7__5_ CARRYB_6__5_ SUMB_6__6_ CARRYB_7__5_ SUMB_7__5_ VDD VSS FA_X1 
XS2_7_4 ab_7__4_ CARRYB_6__4_ SUMB_6__5_ CARRYB_7__4_ SUMB_7__4_ VDD VSS FA_X1 
XS2_7_3 ab_7__3_ CARRYB_6__3_ SUMB_6__4_ CARRYB_7__3_ SUMB_7__3_ VDD VSS FA_X1 
XS2_7_2 ab_7__2_ CARRYB_6__2_ SUMB_6__3_ CARRYB_7__2_ SUMB_7__2_ VDD VSS FA_X1 
XS2_7_1 ab_7__1_ CARRYB_6__1_ SUMB_6__2_ CARRYB_7__1_ SUMB_7__1_ VDD VSS FA_X1 
XS1_7_0 ab_7__0_ CARRYB_6__0_ SUMB_6__1_ CARRYB_7__0_ PRODUCT[7] VDD VSS FA_X1 
XS3_8_16 ab_8__16_ CARRYB_7__16_ ab_7__17_ CARRYB_8__16_ SUMB_8__16_ VDD VSS FA_X1 
XS2_8_15 ab_8__15_ CARRYB_7__15_ SUMB_7__16_ CARRYB_8__15_ SUMB_8__15_ VDD VSS FA_X1 
XS2_8_14 ab_8__14_ CARRYB_7__14_ SUMB_7__15_ CARRYB_8__14_ SUMB_8__14_ VDD VSS FA_X1 
XS2_8_13 ab_8__13_ CARRYB_7__13_ SUMB_7__14_ CARRYB_8__13_ SUMB_8__13_ VDD VSS FA_X1 
XS2_8_12 ab_8__12_ CARRYB_7__12_ SUMB_7__13_ CARRYB_8__12_ SUMB_8__12_ VDD VSS FA_X1 
XS2_8_11 ab_8__11_ CARRYB_7__11_ SUMB_7__12_ CARRYB_8__11_ SUMB_8__11_ VDD VSS FA_X1 
XS2_8_10 ab_8__10_ CARRYB_7__10_ SUMB_7__11_ CARRYB_8__10_ SUMB_8__10_ VDD VSS FA_X1 
XS2_8_9 ab_8__9_ CARRYB_7__9_ SUMB_7__10_ CARRYB_8__9_ SUMB_8__9_ VDD VSS FA_X1 
XS2_8_8 ab_8__8_ CARRYB_7__8_ SUMB_7__9_ CARRYB_8__8_ SUMB_8__8_ VDD VSS FA_X1 
XS2_8_7 ab_8__7_ CARRYB_7__7_ SUMB_7__8_ CARRYB_8__7_ SUMB_8__7_ VDD VSS FA_X1 
XS2_8_6 ab_8__6_ CARRYB_7__6_ SUMB_7__7_ CARRYB_8__6_ SUMB_8__6_ VDD VSS FA_X1 
XS2_8_5 ab_8__5_ CARRYB_7__5_ SUMB_7__6_ CARRYB_8__5_ SUMB_8__5_ VDD VSS FA_X1 
XS2_8_4 ab_8__4_ CARRYB_7__4_ SUMB_7__5_ CARRYB_8__4_ SUMB_8__4_ VDD VSS FA_X1 
XS2_8_3 ab_8__3_ CARRYB_7__3_ SUMB_7__4_ CARRYB_8__3_ SUMB_8__3_ VDD VSS FA_X1 
XS2_8_2 ab_8__2_ CARRYB_7__2_ SUMB_7__3_ CARRYB_8__2_ SUMB_8__2_ VDD VSS FA_X1 
XS2_8_1 ab_8__1_ CARRYB_7__1_ SUMB_7__2_ CARRYB_8__1_ SUMB_8__1_ VDD VSS FA_X1 
XS1_8_0 ab_8__0_ CARRYB_7__0_ SUMB_7__1_ CARRYB_8__0_ PRODUCT[8] VDD VSS FA_X1 
XS3_9_16 ab_9__16_ CARRYB_8__16_ ab_8__17_ CARRYB_9__16_ SUMB_9__16_ VDD VSS FA_X1 
XS2_9_15 ab_9__15_ CARRYB_8__15_ SUMB_8__16_ CARRYB_9__15_ SUMB_9__15_ VDD VSS FA_X1 
XS2_9_14 ab_9__14_ CARRYB_8__14_ SUMB_8__15_ CARRYB_9__14_ SUMB_9__14_ VDD VSS FA_X1 
XS2_9_13 ab_9__13_ CARRYB_8__13_ SUMB_8__14_ CARRYB_9__13_ SUMB_9__13_ VDD VSS FA_X1 
XS2_9_12 ab_9__12_ CARRYB_8__12_ SUMB_8__13_ CARRYB_9__12_ SUMB_9__12_ VDD VSS FA_X1 
XU63 CARRYB_15__5_ SUMB_15__6_ n62 VDD VSS XOR2_X1 
XU62 CARRYB_15__15_ SUMB_15__16_ n61 VDD VSS AND2_X1 
XU61 CARRYB_15__14_ SUMB_15__15_ n60 VDD VSS AND2_X1 
XU60 CARRYB_15__13_ SUMB_15__14_ n59 VDD VSS AND2_X1 
XU59 CARRYB_15__12_ SUMB_15__13_ n58 VDD VSS AND2_X1 
XU58 CARRYB_15__11_ SUMB_15__12_ n57 VDD VSS AND2_X1 
XU57 CARRYB_15__10_ SUMB_15__11_ n56 VDD VSS AND2_X1 
XU56 CARRYB_15__9_ SUMB_15__10_ n55 VDD VSS AND2_X1 
XU55 CARRYB_15__8_ SUMB_15__9_ n54 VDD VSS AND2_X1 
XU54 CARRYB_15__7_ SUMB_15__8_ n53 VDD VSS AND2_X1 
XU53 CARRYB_15__6_ SUMB_15__7_ n52 VDD VSS AND2_X1 
XU52 CARRYB_15__5_ SUMB_15__6_ n51 VDD VSS AND2_X1 
XU51 CARRYB_15__4_ SUMB_15__5_ n50 VDD VSS AND2_X1 
XU50 CARRYB_15__16_ SUMB_15__17_ n49 VDD VSS AND2_X1 
XU49 CARRYB_15__16_ SUMB_15__17_ n48 VDD VSS XOR2_X1 
XU48 CARRYB_15__14_ SUMB_15__15_ n47 VDD VSS XOR2_X1 
XU47 CARRYB_15__12_ SUMB_15__13_ n46 VDD VSS XOR2_X1 
XU46 CARRYB_15__10_ SUMB_15__11_ n45 VDD VSS XOR2_X1 
XU45 CARRYB_15__8_ SUMB_15__9_ n44 VDD VSS XOR2_X1 
XU44 CARRYB_15__6_ SUMB_15__7_ n43 VDD VSS XOR2_X1 
XU43 CARRYB_15__3_ SUMB_15__4_ n42 VDD VSS XOR2_X1 
XU42 CARRYB_15__3_ SUMB_15__4_ n41 VDD VSS AND2_X1 
XU41 CARRYB_15__2_ SUMB_15__3_ n40 VDD VSS AND2_X1 
XU40 CARRYB_15__0_ SUMB_15__1_ n39 VDD VSS AND2_X1 
XU39 CARRYB_15__0_ SUMB_15__1_ n38 VDD VSS XOR2_X1 
XU38 CARRYB_15__4_ SUMB_15__5_ n37 VDD VSS XOR2_X1 
XU37 CARRYB_15__2_ SUMB_15__3_ n36 VDD VSS XOR2_X1 
XU36 ab_1__0_ ab_0__1_ PRODUCT[1] VDD VSS XOR2_X1 
XU35 CARRYB_15__17_ n70 VDD VSS INV_X1 
XU34 ab_1__1_ ab_0__2_ n34 VDD VSS XOR2_X1 
XU33 ab_1__2_ ab_0__3_ n33 VDD VSS XOR2_X1 
XU32 ab_1__16_ ab_0__17_ n32 VDD VSS XOR2_X1 
XU31 ab_1__3_ ab_0__4_ n31 VDD VSS XOR2_X1 
XU30 ab_1__4_ ab_0__5_ n30 VDD VSS XOR2_X1 
XU29 ab_1__5_ ab_0__6_ n29 VDD VSS XOR2_X1 
XU28 ab_1__6_ ab_0__7_ n28 VDD VSS XOR2_X1 
XU27 ab_1__7_ ab_0__8_ n27 VDD VSS XOR2_X1 
XU26 ab_1__8_ ab_0__9_ n26 VDD VSS XOR2_X1 
XU25 ab_1__9_ ab_0__10_ n25 VDD VSS XOR2_X1 
XU24 ab_1__10_ ab_0__11_ n24 VDD VSS XOR2_X1 
XU23 ab_1__11_ ab_0__12_ n23 VDD VSS XOR2_X1 
XU22 ab_1__12_ ab_0__13_ n22 VDD VSS XOR2_X1 
XU21 ab_1__13_ ab_0__14_ n21 VDD VSS XOR2_X1 
XU20 ab_1__14_ ab_0__15_ n20 VDD VSS XOR2_X1 
XU19 ab_1__15_ ab_0__16_ n19 VDD VSS XOR2_X1 
XU18 ab_0__17_ ab_1__16_ n18 VDD VSS AND2_X1 
XU17 ab_0__1_ ab_1__0_ n17 VDD VSS AND2_X1 
XU16 ab_0__2_ ab_1__1_ n16 VDD VSS AND2_X1 
XU15 ab_0__3_ ab_1__2_ n15 VDD VSS AND2_X1 
XU14 ab_0__4_ ab_1__3_ n14 VDD VSS AND2_X1 
XU13 ab_0__5_ ab_1__4_ n13 VDD VSS AND2_X1 
XU12 ab_0__6_ ab_1__5_ n12 VDD VSS AND2_X1 
XU11 ab_0__7_ ab_1__6_ n11 VDD VSS AND2_X1 
XU10 ab_0__8_ ab_1__7_ n10 VDD VSS AND2_X1 
XU9 ab_0__9_ ab_1__8_ n9 VDD VSS AND2_X1 
XU8 ab_0__10_ ab_1__9_ n8 VDD VSS AND2_X1 
XU7 ab_0__11_ ab_1__10_ n7 VDD VSS AND2_X1 
XU6 ab_0__12_ ab_1__11_ n6 VDD VSS AND2_X1 
XU5 ab_0__13_ ab_1__12_ n5 VDD VSS AND2_X1 
XU4 ab_0__14_ ab_1__13_ n4 VDD VSS AND2_X1 
XU3 ab_0__15_ ab_1__14_ n3 VDD VSS AND2_X1 
XU2 ab_0__16_ ab_1__15_ n2 VDD VSS AND2_X1 
XS3_2_16 ab_2__16_ n18 ab_1__17_ CARRYB_2__16_ SUMB_2__16_ VDD VSS FA_X1 
XS2_2_15 ab_2__15_ n2 n32 CARRYB_2__15_ SUMB_2__15_ VDD VSS FA_X1 
XS2_2_14 ab_2__14_ n3 n19 CARRYB_2__14_ SUMB_2__14_ VDD VSS FA_X1 
XS2_2_13 ab_2__13_ n4 n20 CARRYB_2__13_ SUMB_2__13_ VDD VSS FA_X1 
XS2_2_12 ab_2__12_ n5 n21 CARRYB_2__12_ SUMB_2__12_ VDD VSS FA_X1 
XS2_2_11 ab_2__11_ n6 n22 CARRYB_2__11_ SUMB_2__11_ VDD VSS FA_X1 
XS2_2_10 ab_2__10_ n7 n23 CARRYB_2__10_ SUMB_2__10_ VDD VSS FA_X1 
XS2_2_9 ab_2__9_ n8 n24 CARRYB_2__9_ SUMB_2__9_ VDD VSS FA_X1 
XS2_2_8 ab_2__8_ n9 n25 CARRYB_2__8_ SUMB_2__8_ VDD VSS FA_X1 
XS2_2_7 ab_2__7_ n10 n26 CARRYB_2__7_ SUMB_2__7_ VDD VSS FA_X1 
XS2_2_6 ab_2__6_ n11 n27 CARRYB_2__6_ SUMB_2__6_ VDD VSS FA_X1 
XS2_2_5 ab_2__5_ n12 n28 CARRYB_2__5_ SUMB_2__5_ VDD VSS FA_X1 
XS2_2_4 ab_2__4_ n13 n29 CARRYB_2__4_ SUMB_2__4_ VDD VSS FA_X1 
XS2_2_3 ab_2__3_ n14 n30 CARRYB_2__3_ SUMB_2__3_ VDD VSS FA_X1 
XS2_2_2 ab_2__2_ n15 n31 CARRYB_2__2_ SUMB_2__2_ VDD VSS FA_X1 
XS2_2_1 ab_2__1_ n16 n33 CARRYB_2__1_ SUMB_2__1_ VDD VSS FA_X1 
XS1_2_0 ab_2__0_ n17 n34 CARRYB_2__0_ PRODUCT[2] VDD VSS FA_X1 
XS3_3_16 ab_3__16_ CARRYB_2__16_ ab_2__17_ CARRYB_3__16_ SUMB_3__16_ VDD VSS FA_X1 
XS2_3_15 ab_3__15_ CARRYB_2__15_ SUMB_2__16_ CARRYB_3__15_ SUMB_3__15_ VDD VSS FA_X1 
XS2_3_14 ab_3__14_ CARRYB_2__14_ SUMB_2__15_ CARRYB_3__14_ SUMB_3__14_ VDD VSS FA_X1 
XS2_3_13 ab_3__13_ CARRYB_2__13_ SUMB_2__14_ CARRYB_3__13_ SUMB_3__13_ VDD VSS FA_X1 
XS2_3_12 ab_3__12_ CARRYB_2__12_ SUMB_2__13_ CARRYB_3__12_ SUMB_3__12_ VDD VSS FA_X1 
XS2_3_11 ab_3__11_ CARRYB_2__11_ SUMB_2__12_ CARRYB_3__11_ SUMB_3__11_ VDD VSS FA_X1 
XS2_3_10 ab_3__10_ CARRYB_2__10_ SUMB_2__11_ CARRYB_3__10_ SUMB_3__10_ VDD VSS FA_X1 
XS2_3_9 ab_3__9_ CARRYB_2__9_ SUMB_2__10_ CARRYB_3__9_ SUMB_3__9_ VDD VSS FA_X1 
XS2_3_8 ab_3__8_ CARRYB_2__8_ SUMB_2__9_ CARRYB_3__8_ SUMB_3__8_ VDD VSS FA_X1 
XS2_3_7 ab_3__7_ CARRYB_2__7_ SUMB_2__8_ CARRYB_3__7_ SUMB_3__7_ VDD VSS FA_X1 
XS2_3_6 ab_3__6_ CARRYB_2__6_ SUMB_2__7_ CARRYB_3__6_ SUMB_3__6_ VDD VSS FA_X1 
XS2_3_5 ab_3__5_ CARRYB_2__5_ SUMB_2__6_ CARRYB_3__5_ SUMB_3__5_ VDD VSS FA_X1 
XS2_3_4 ab_3__4_ CARRYB_2__4_ SUMB_2__5_ CARRYB_3__4_ SUMB_3__4_ VDD VSS FA_X1 
XS2_3_3 ab_3__3_ CARRYB_2__3_ SUMB_2__4_ CARRYB_3__3_ SUMB_3__3_ VDD VSS FA_X1 
XU156 n91 n77 ab_7__11_ VDD VSS NOR2_X1 
XU155 n90 n77 ab_7__12_ VDD VSS NOR2_X1 
XU154 n89 n77 ab_7__13_ VDD VSS NOR2_X1 
XU153 n88 n77 ab_7__14_ VDD VSS NOR2_X1 
XU152 n87 n77 ab_7__15_ VDD VSS NOR2_X1 
XU151 n86 n77 ab_7__16_ VDD VSS NOR2_X1 
XU150 A[7] n85 ab_7__17_ VDD VSS NOR2_X1 
XU149 n101 n77 ab_7__1_ VDD VSS NOR2_X1 
XU148 n100 n77 ab_7__2_ VDD VSS NOR2_X1 
XU147 n99 n77 ab_7__3_ VDD VSS NOR2_X1 
XU146 n98 n77 ab_7__4_ VDD VSS NOR2_X1 
XU145 n97 n77 ab_7__5_ VDD VSS NOR2_X1 
XU144 n96 n77 ab_7__6_ VDD VSS NOR2_X1 
XU143 n95 n77 ab_7__7_ VDD VSS NOR2_X1 
XU142 n94 n77 ab_7__8_ VDD VSS NOR2_X1 
XU141 n93 n77 ab_7__9_ VDD VSS NOR2_X1 
XU140 n102 n76 ab_8__0_ VDD VSS NOR2_X1 
XU139 n92 n76 ab_8__10_ VDD VSS NOR2_X1 
XU138 n91 n76 ab_8__11_ VDD VSS NOR2_X1 
XU137 n90 n76 ab_8__12_ VDD VSS NOR2_X1 
XU136 n89 n76 ab_8__13_ VDD VSS NOR2_X1 
XU135 n88 n76 ab_8__14_ VDD VSS NOR2_X1 
XU134 n87 n76 ab_8__15_ VDD VSS NOR2_X1 
XU133 n86 n76 ab_8__16_ VDD VSS NOR2_X1 
XU132 A[8] n85 ab_8__17_ VDD VSS NOR2_X1 
XU131 n101 n76 ab_8__1_ VDD VSS NOR2_X1 
XU130 n100 n76 ab_8__2_ VDD VSS NOR2_X1 
XU129 n99 n76 ab_8__3_ VDD VSS NOR2_X1 
XU128 n98 n76 ab_8__4_ VDD VSS NOR2_X1 
XU127 n97 n76 ab_8__5_ VDD VSS NOR2_X1 
XU126 n96 n76 ab_8__6_ VDD VSS NOR2_X1 
XU125 n95 n76 ab_8__7_ VDD VSS NOR2_X1 
XU124 n94 n76 ab_8__8_ VDD VSS NOR2_X1 
XU123 n93 n76 ab_8__9_ VDD VSS NOR2_X1 
XU122 n75 n102 ab_9__0_ VDD VSS NOR2_X1 
XU121 n75 n92 ab_9__10_ VDD VSS NOR2_X1 
XU120 n75 n91 ab_9__11_ VDD VSS NOR2_X1 
XU119 n75 n90 ab_9__12_ VDD VSS NOR2_X1 
XU118 n75 n89 ab_9__13_ VDD VSS NOR2_X1 
XU117 n75 n88 ab_9__14_ VDD VSS NOR2_X1 
XU116 n75 n87 ab_9__15_ VDD VSS NOR2_X1 
XU115 n75 n86 ab_9__16_ VDD VSS NOR2_X1 
XU114 A[9] n85 ab_9__17_ VDD VSS NOR2_X1 
XU113 n75 n101 ab_9__1_ VDD VSS NOR2_X1 
XU112 n75 n100 ab_9__2_ VDD VSS NOR2_X1 
XU111 n75 n99 ab_9__3_ VDD VSS NOR2_X1 
XU110 n75 n98 ab_9__4_ VDD VSS NOR2_X1 
XU109 n75 n97 ab_9__5_ VDD VSS NOR2_X1 
XU108 n75 n96 ab_9__6_ VDD VSS NOR2_X1 
XU107 n75 n95 ab_9__7_ VDD VSS NOR2_X1 
XU106 n75 n94 ab_9__8_ VDD VSS NOR2_X1 
XU105 n75 n93 ab_9__9_ VDD VSS NOR2_X1 
XU101 A[15] SUMB_15__0_ PRODUCT[15] VDD VSS XOR2_X1 
XU89 A[15] SUMB_15__0_ n68 VDD VSS AND2_X1 
XU68 CARRYB_15__15_ SUMB_15__16_ n67 VDD VSS XOR2_X1 
XU67 CARRYB_15__13_ SUMB_15__14_ n66 VDD VSS XOR2_X1 
XU66 CARRYB_15__11_ SUMB_15__12_ n65 VDD VSS XOR2_X1 
XU65 CARRYB_15__9_ SUMB_15__10_ n64 VDD VSS XOR2_X1 
XU64 CARRYB_15__7_ SUMB_15__8_ n63 VDD VSS XOR2_X1 
XU249 n93 n83 ab_1__9_ VDD VSS NOR2_X1 
XU248 n102 n82 ab_2__0_ VDD VSS NOR2_X1 
XU247 n92 n82 ab_2__10_ VDD VSS NOR2_X1 
XU246 n91 n82 ab_2__11_ VDD VSS NOR2_X1 
XU245 n90 n82 ab_2__12_ VDD VSS NOR2_X1 
XU244 n89 n82 ab_2__13_ VDD VSS NOR2_X1 
XU243 n88 n82 ab_2__14_ VDD VSS NOR2_X1 
XU242 n87 n82 ab_2__15_ VDD VSS NOR2_X1 
XU241 n86 n82 ab_2__16_ VDD VSS NOR2_X1 
XU240 A[2] n85 ab_2__17_ VDD VSS NOR2_X1 
XU239 n101 n82 ab_2__1_ VDD VSS NOR2_X1 
XU238 n100 n82 ab_2__2_ VDD VSS NOR2_X1 
XU237 n99 n82 ab_2__3_ VDD VSS NOR2_X1 
XU236 n98 n82 ab_2__4_ VDD VSS NOR2_X1 
XU235 n97 n82 ab_2__5_ VDD VSS NOR2_X1 
XU234 n96 n82 ab_2__6_ VDD VSS NOR2_X1 
XU233 n95 n82 ab_2__7_ VDD VSS NOR2_X1 
XU232 n94 n82 ab_2__8_ VDD VSS NOR2_X1 
XU231 n93 n82 ab_2__9_ VDD VSS NOR2_X1 
XU230 n102 n81 ab_3__0_ VDD VSS NOR2_X1 
XU229 n92 n81 ab_3__10_ VDD VSS NOR2_X1 
XU228 n91 n81 ab_3__11_ VDD VSS NOR2_X1 
XU227 n90 n81 ab_3__12_ VDD VSS NOR2_X1 
XU226 n89 n81 ab_3__13_ VDD VSS NOR2_X1 
XU225 n88 n81 ab_3__14_ VDD VSS NOR2_X1 
XU224 n87 n81 ab_3__15_ VDD VSS NOR2_X1 
XU223 n86 n81 ab_3__16_ VDD VSS NOR2_X1 
XU222 A[3] n85 ab_3__17_ VDD VSS NOR2_X1 
XU221 n101 n81 ab_3__1_ VDD VSS NOR2_X1 
XU220 n100 n81 ab_3__2_ VDD VSS NOR2_X1 
XU219 n99 n81 ab_3__3_ VDD VSS NOR2_X1 
XU218 n98 n81 ab_3__4_ VDD VSS NOR2_X1 
XU217 n97 n81 ab_3__5_ VDD VSS NOR2_X1 
XU216 n96 n81 ab_3__6_ VDD VSS NOR2_X1 
XU215 n95 n81 ab_3__7_ VDD VSS NOR2_X1 
XU214 n94 n81 ab_3__8_ VDD VSS NOR2_X1 
XU213 n93 n81 ab_3__9_ VDD VSS NOR2_X1 
XU212 n102 n80 ab_4__0_ VDD VSS NOR2_X1 
XU211 n92 n80 ab_4__10_ VDD VSS NOR2_X1 
XU210 n91 n80 ab_4__11_ VDD VSS NOR2_X1 
XU209 n90 n80 ab_4__12_ VDD VSS NOR2_X1 
XU208 n89 n80 ab_4__13_ VDD VSS NOR2_X1 
XU207 n88 n80 ab_4__14_ VDD VSS NOR2_X1 
XU206 n87 n80 ab_4__15_ VDD VSS NOR2_X1 
XU205 n86 n80 ab_4__16_ VDD VSS NOR2_X1 
XU204 A[4] n85 ab_4__17_ VDD VSS NOR2_X1 
XU203 n101 n80 ab_4__1_ VDD VSS NOR2_X1 
XU202 n100 n80 ab_4__2_ VDD VSS NOR2_X1 
XU201 n99 n80 ab_4__3_ VDD VSS NOR2_X1 
XU200 n98 n80 ab_4__4_ VDD VSS NOR2_X1 
XU199 n97 n80 ab_4__5_ VDD VSS NOR2_X1 
XU198 n96 n80 ab_4__6_ VDD VSS NOR2_X1 
XU197 n95 n80 ab_4__7_ VDD VSS NOR2_X1 
XU196 n94 n80 ab_4__8_ VDD VSS NOR2_X1 
XU195 n93 n80 ab_4__9_ VDD VSS NOR2_X1 
XU194 n102 n79 ab_5__0_ VDD VSS NOR2_X1 
XU193 n92 n79 ab_5__10_ VDD VSS NOR2_X1 
XU192 n91 n79 ab_5__11_ VDD VSS NOR2_X1 
XU191 n90 n79 ab_5__12_ VDD VSS NOR2_X1 
XU190 n89 n79 ab_5__13_ VDD VSS NOR2_X1 
XU189 n88 n79 ab_5__14_ VDD VSS NOR2_X1 
XU188 n87 n79 ab_5__15_ VDD VSS NOR2_X1 
XU187 n86 n79 ab_5__16_ VDD VSS NOR2_X1 
XU186 A[5] n85 ab_5__17_ VDD VSS NOR2_X1 
XU185 n101 n79 ab_5__1_ VDD VSS NOR2_X1 
XU184 n100 n79 ab_5__2_ VDD VSS NOR2_X1 
XU183 n99 n79 ab_5__3_ VDD VSS NOR2_X1 
XU182 n98 n79 ab_5__4_ VDD VSS NOR2_X1 
XU181 n97 n79 ab_5__5_ VDD VSS NOR2_X1 
XU180 n96 n79 ab_5__6_ VDD VSS NOR2_X1 
XU179 n95 n79 ab_5__7_ VDD VSS NOR2_X1 
XU178 n94 n79 ab_5__8_ VDD VSS NOR2_X1 
XU177 n93 n79 ab_5__9_ VDD VSS NOR2_X1 
XU176 n102 n78 ab_6__0_ VDD VSS NOR2_X1 
XU175 n92 n78 ab_6__10_ VDD VSS NOR2_X1 
XU174 n91 n78 ab_6__11_ VDD VSS NOR2_X1 
XU173 n90 n78 ab_6__12_ VDD VSS NOR2_X1 
XU172 n89 n78 ab_6__13_ VDD VSS NOR2_X1 
XU171 n88 n78 ab_6__14_ VDD VSS NOR2_X1 
XU170 n87 n78 ab_6__15_ VDD VSS NOR2_X1 
XU169 n86 n78 ab_6__16_ VDD VSS NOR2_X1 
XU168 A[6] n85 ab_6__17_ VDD VSS NOR2_X1 
XU167 n101 n78 ab_6__1_ VDD VSS NOR2_X1 
XU166 n100 n78 ab_6__2_ VDD VSS NOR2_X1 
XU165 n99 n78 ab_6__3_ VDD VSS NOR2_X1 
XU164 n98 n78 ab_6__4_ VDD VSS NOR2_X1 
XU163 n97 n78 ab_6__5_ VDD VSS NOR2_X1 
XU162 n96 n78 ab_6__6_ VDD VSS NOR2_X1 
XU161 n95 n78 ab_6__7_ VDD VSS NOR2_X1 
XU160 n94 n78 ab_6__8_ VDD VSS NOR2_X1 
XU159 n93 n78 ab_6__9_ VDD VSS NOR2_X1 
XU158 n102 n77 ab_7__0_ VDD VSS NOR2_X1 
XU157 n92 n77 ab_7__10_ VDD VSS NOR2_X1 
XU342 n96 n73 ab_11__6_ VDD VSS NOR2_X1 
XU341 n95 n73 ab_11__7_ VDD VSS NOR2_X1 
XU340 n94 n73 ab_11__8_ VDD VSS NOR2_X1 
XU339 n93 n73 ab_11__9_ VDD VSS NOR2_X1 
XU338 n102 n72 ab_12__0_ VDD VSS NOR2_X1 
XU337 n92 n72 ab_12__10_ VDD VSS NOR2_X1 
XU336 n91 n72 ab_12__11_ VDD VSS NOR2_X1 
XU335 n90 n72 ab_12__12_ VDD VSS NOR2_X1 
XU334 n89 n72 ab_12__13_ VDD VSS NOR2_X1 
XU333 n88 n72 ab_12__14_ VDD VSS NOR2_X1 
XU332 n87 n72 ab_12__15_ VDD VSS NOR2_X1 
XU331 n86 n72 ab_12__16_ VDD VSS NOR2_X1 
XU330 A[12] n85 ab_12__17_ VDD VSS NOR2_X1 
XU329 n101 n72 ab_12__1_ VDD VSS NOR2_X1 
XU328 n100 n72 ab_12__2_ VDD VSS NOR2_X1 
XU327 n99 n72 ab_12__3_ VDD VSS NOR2_X1 
XU326 n98 n72 ab_12__4_ VDD VSS NOR2_X1 
XU325 n97 n72 ab_12__5_ VDD VSS NOR2_X1 
XU324 n96 n72 ab_12__6_ VDD VSS NOR2_X1 
XU323 n95 n72 ab_12__7_ VDD VSS NOR2_X1 
XU322 n94 n72 ab_12__8_ VDD VSS NOR2_X1 
XU321 n93 n72 ab_12__9_ VDD VSS NOR2_X1 
XU320 n102 n71 ab_13__0_ VDD VSS NOR2_X1 
XU319 n92 n71 ab_13__10_ VDD VSS NOR2_X1 
XU318 n91 n71 ab_13__11_ VDD VSS NOR2_X1 
XU317 n90 n71 ab_13__12_ VDD VSS NOR2_X1 
XU316 n89 n71 ab_13__13_ VDD VSS NOR2_X1 
XU315 n88 n71 ab_13__14_ VDD VSS NOR2_X1 
XU314 n87 n71 ab_13__15_ VDD VSS NOR2_X1 
XU313 n86 n71 ab_13__16_ VDD VSS NOR2_X1 
XU312 A[13] n85 ab_13__17_ VDD VSS NOR2_X1 
XU311 n101 n71 ab_13__1_ VDD VSS NOR2_X1 
XU310 n100 n71 ab_13__2_ VDD VSS NOR2_X1 
XU309 n99 n71 ab_13__3_ VDD VSS NOR2_X1 
XU308 n98 n71 ab_13__4_ VDD VSS NOR2_X1 
XU307 n97 n71 ab_13__5_ VDD VSS NOR2_X1 
XU306 n96 n71 ab_13__6_ VDD VSS NOR2_X1 
XU305 n95 n71 ab_13__7_ VDD VSS NOR2_X1 
XU304 n94 n71 ab_13__8_ VDD VSS NOR2_X1 
XU303 n93 n71 ab_13__9_ VDD VSS NOR2_X1 
XU302 n102 n35 ab_14__0_ VDD VSS NOR2_X1 
XU301 n92 n35 ab_14__10_ VDD VSS NOR2_X1 
XU300 n91 n35 ab_14__11_ VDD VSS NOR2_X1 
XU299 n90 n35 ab_14__12_ VDD VSS NOR2_X1 
XU298 n89 n35 ab_14__13_ VDD VSS NOR2_X1 
XU297 n88 n35 ab_14__14_ VDD VSS NOR2_X1 
XU296 n87 n35 ab_14__15_ VDD VSS NOR2_X1 
XU295 n86 n35 ab_14__16_ VDD VSS NOR2_X1 
XU294 A[14] n85 ab_14__17_ VDD VSS NOR2_X1 
XU293 n101 n35 ab_14__1_ VDD VSS NOR2_X1 
XU292 n100 n35 ab_14__2_ VDD VSS NOR2_X1 
XU291 n99 n35 ab_14__3_ VDD VSS NOR2_X1 
XU290 n98 n35 ab_14__4_ VDD VSS NOR2_X1 
XU289 n97 n35 ab_14__5_ VDD VSS NOR2_X1 
XU288 n96 n35 ab_14__6_ VDD VSS NOR2_X1 
XU287 n95 n35 ab_14__7_ VDD VSS NOR2_X1 
XU286 n94 n35 ab_14__8_ VDD VSS NOR2_X1 
XU285 n93 n35 ab_14__9_ VDD VSS NOR2_X1 
XU284 B[0] n1 ab_15__0_ VDD VSS NOR2_X1 
XU283 B[10] n1 ab_15__10_ VDD VSS NOR2_X1 
XU282 B[11] n1 ab_15__11_ VDD VSS NOR2_X1 
XU281 B[12] n1 ab_15__12_ VDD VSS NOR2_X1 
XU280 B[13] n1 ab_15__13_ VDD VSS NOR2_X1 
XU279 B[14] n1 ab_15__14_ VDD VSS NOR2_X1 
XU278 B[15] n1 ab_15__15_ VDD VSS NOR2_X1 
XU277 B[16] n1 ab_15__16_ VDD VSS NOR2_X1 
XU276 n85 n1 ab_15__17_ VDD VSS NOR2_X1 
XU275 B[1] n1 ab_15__1_ VDD VSS NOR2_X1 
XU274 B[2] n1 ab_15__2_ VDD VSS NOR2_X1 
XU273 B[3] n1 ab_15__3_ VDD VSS NOR2_X1 
XU272 B[4] n1 ab_15__4_ VDD VSS NOR2_X1 
XU271 B[5] n1 ab_15__5_ VDD VSS NOR2_X1 
XU270 B[6] n1 ab_15__6_ VDD VSS NOR2_X1 
XU269 B[7] n1 ab_15__7_ VDD VSS NOR2_X1 
XU268 B[8] n1 ab_15__8_ VDD VSS NOR2_X1 
XU267 B[9] n1 ab_15__9_ VDD VSS NOR2_X1 
XU266 n102 n83 ab_1__0_ VDD VSS NOR2_X1 
XU265 n92 n83 ab_1__10_ VDD VSS NOR2_X1 
XU264 n91 n83 ab_1__11_ VDD VSS NOR2_X1 
XU263 n90 n83 ab_1__12_ VDD VSS NOR2_X1 
XU262 n89 n83 ab_1__13_ VDD VSS NOR2_X1 
XU261 n88 n83 ab_1__14_ VDD VSS NOR2_X1 
XU260 n87 n83 ab_1__15_ VDD VSS NOR2_X1 
XU259 n86 n83 ab_1__16_ VDD VSS NOR2_X1 
XU258 A[1] n85 ab_1__17_ VDD VSS NOR2_X1 
XU257 n101 n83 ab_1__1_ VDD VSS NOR2_X1 
XU256 n100 n83 ab_1__2_ VDD VSS NOR2_X1 
XU255 n99 n83 ab_1__3_ VDD VSS NOR2_X1 
XU254 n98 n83 ab_1__4_ VDD VSS NOR2_X1 
XU253 n97 n83 ab_1__5_ VDD VSS NOR2_X1 
XU252 n96 n83 ab_1__6_ VDD VSS NOR2_X1 
XU251 n95 n83 ab_1__7_ VDD VSS NOR2_X1 
XU250 n94 n83 ab_1__8_ VDD VSS NOR2_X1 
XU392 n102 n84 PRODUCT[0] VDD VSS NOR2_X1 
XU391 n92 n84 ab_0__10_ VDD VSS NOR2_X1 
XU390 n91 n84 ab_0__11_ VDD VSS NOR2_X1 
XU389 n90 n84 ab_0__12_ VDD VSS NOR2_X1 
XU388 n89 n84 ab_0__13_ VDD VSS NOR2_X1 
XU387 n88 n84 ab_0__14_ VDD VSS NOR2_X1 
XU386 n87 n84 ab_0__15_ VDD VSS NOR2_X1 
XU385 n86 n84 ab_0__16_ VDD VSS NOR2_X1 
XU384 A[0] n85 ab_0__17_ VDD VSS NOR2_X1 
XU383 n101 n84 ab_0__1_ VDD VSS NOR2_X1 
XU382 n100 n84 ab_0__2_ VDD VSS NOR2_X1 
XU381 n99 n84 ab_0__3_ VDD VSS NOR2_X1 
XU380 n98 n84 ab_0__4_ VDD VSS NOR2_X1 
XU379 n97 n84 ab_0__5_ VDD VSS NOR2_X1 
XU378 n96 n84 ab_0__6_ VDD VSS NOR2_X1 
XU377 n95 n84 ab_0__7_ VDD VSS NOR2_X1 
XU376 n94 n84 ab_0__8_ VDD VSS NOR2_X1 
XU375 n93 n84 ab_0__9_ VDD VSS NOR2_X1 
XU374 n102 n74 ab_10__0_ VDD VSS NOR2_X1 
XU373 n92 n74 ab_10__10_ VDD VSS NOR2_X1 
XU372 n91 n74 ab_10__11_ VDD VSS NOR2_X1 
XU371 n90 n74 ab_10__12_ VDD VSS NOR2_X1 
XU370 n89 n74 ab_10__13_ VDD VSS NOR2_X1 
XU369 n88 n74 ab_10__14_ VDD VSS NOR2_X1 
XU368 n87 n74 ab_10__15_ VDD VSS NOR2_X1 
XU367 n86 n74 ab_10__16_ VDD VSS NOR2_X1 
XU366 A[10] n85 ab_10__17_ VDD VSS NOR2_X1 
XU365 n101 n74 ab_10__1_ VDD VSS NOR2_X1 
XU364 n100 n74 ab_10__2_ VDD VSS NOR2_X1 
XU363 n99 n74 ab_10__3_ VDD VSS NOR2_X1 
XU362 n98 n74 ab_10__4_ VDD VSS NOR2_X1 
XU361 n97 n74 ab_10__5_ VDD VSS NOR2_X1 
XU360 n96 n74 ab_10__6_ VDD VSS NOR2_X1 
XU359 n95 n74 ab_10__7_ VDD VSS NOR2_X1 
XU358 n94 n74 ab_10__8_ VDD VSS NOR2_X1 
XU357 n93 n74 ab_10__9_ VDD VSS NOR2_X1 
XU356 n102 n73 ab_11__0_ VDD VSS NOR2_X1 
XU355 n92 n73 ab_11__10_ VDD VSS NOR2_X1 
XU354 n91 n73 ab_11__11_ VDD VSS NOR2_X1 
XU353 n90 n73 ab_11__12_ VDD VSS NOR2_X1 
XU352 n89 n73 ab_11__13_ VDD VSS NOR2_X1 
XU351 n88 n73 ab_11__14_ VDD VSS NOR2_X1 
XU350 n87 n73 ab_11__15_ VDD VSS NOR2_X1 
XU349 n86 n73 ab_11__16_ VDD VSS NOR2_X1 
XU348 A[11] n85 ab_11__17_ VDD VSS NOR2_X1 
XU347 n101 n73 ab_11__1_ VDD VSS NOR2_X1 
XU346 n100 n73 ab_11__2_ VDD VSS NOR2_X1 
XU345 n99 n73 ab_11__3_ VDD VSS NOR2_X1 
XU344 n98 n73 ab_11__4_ VDD VSS NOR2_X1 
XU343 n97 n73 ab_11__5_ VDD VSS NOR2_X1 
XU1 A[15] n1 VDD VSS INV_X1 
XU69 A[14] n35 VDD VSS INV_X1 
XU70 A[13] n71 VDD VSS INV_X1 
XU71 A[12] n72 VDD VSS INV_X1 
XU72 A[11] n73 VDD VSS INV_X1 
XU73 A[10] n74 VDD VSS INV_X1 
XU74 A[9] n75 VDD VSS INV_X1 
XU75 A[8] n76 VDD VSS INV_X1 
XU76 A[7] n77 VDD VSS INV_X1 
XU77 A[6] n78 VDD VSS INV_X1 
XU78 A[5] n79 VDD VSS INV_X1 
XU79 A[4] n80 VDD VSS INV_X1 
XU80 A[3] n81 VDD VSS INV_X1 
XU81 A[2] n82 VDD VSS INV_X1 
XU82 A[1] n83 VDD VSS INV_X1 
XU83 A[0] n84 VDD VSS INV_X1 
XU84 B[17] n85 VDD VSS INV_X1 
XU85 B[16] n86 VDD VSS INV_X1 
XU86 B[15] n87 VDD VSS INV_X1 
XU87 B[14] n88 VDD VSS INV_X1 
XU88 B[13] n89 VDD VSS INV_X1 
XU90 B[12] n90 VDD VSS INV_X1 
XU91 B[11] n91 VDD VSS INV_X1 
XU92 B[10] n92 VDD VSS INV_X1 
XU93 B[9] n93 VDD VSS INV_X1 
XU94 B[8] n94 VDD VSS INV_X1 
XU95 B[7] n95 VDD VSS INV_X1 
XU96 B[6] n96 VDD VSS INV_X1 
XU97 B[5] n97 VDD VSS INV_X1 
XU98 B[4] n98 VDD VSS INV_X1 
XU99 B[3] n99 VDD VSS INV_X1 
XU100 B[2] n100 VDD VSS INV_X1 
XU102 B[1] n101 VDD VSS INV_X1 
XU103 B[0] n102 VDD VSS INV_X1 
XFS_1 VSS SYNOPSYS_UNCONNECTED_45 VDD VSS PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ n49 n61 n60 n59 n58 n57 n56 n55 n54 n53 n52 n51 n50 n41 n40 A2_16_ n39 n68 VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS n70 n48 n67 n47 n66 n46 n65 
+ n45 n64 n44 n63 n43 n62 n37 n42 n36 A1_15_ n38 PRODUCT[15] PRODUCT[14] PRODUCT[13] 
+ PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] PRODUCT[8] PRODUCT[7] PRODUCT[6] 
+ PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] gng_smul_16_18_DW01_add_0 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37_DW02_mult_0 PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ PRODUCT[15] PRODUCT[14] PRODUCT[13] PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] 
+ PRODUCT[8] PRODUCT[7] PRODUCT[6] PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] PRODUCT[1] 
+ PRODUCT[0] TC VDD VSS B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] 
+ B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] 
+ A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
XU1 A[15] n1 VDD VSS INV_X1 
XS2_11_8 ab_11__8_ CARRYB_10__8_ SUMB_10__9_ CARRYB_11__8_ SUMB_11__8_ VDD VSS FA_X1 
XS2_11_7 ab_11__7_ CARRYB_10__7_ SUMB_10__8_ CARRYB_11__7_ SUMB_11__7_ VDD VSS FA_X1 
XS2_11_6 ab_11__6_ CARRYB_10__6_ SUMB_10__7_ CARRYB_11__6_ SUMB_11__6_ VDD VSS FA_X1 
XS2_11_5 ab_11__5_ CARRYB_10__5_ SUMB_10__6_ CARRYB_11__5_ SUMB_11__5_ VDD VSS FA_X1 
XS2_11_4 ab_11__4_ CARRYB_10__4_ SUMB_10__5_ CARRYB_11__4_ SUMB_11__4_ VDD VSS FA_X1 
XS2_11_3 ab_11__3_ CARRYB_10__3_ SUMB_10__4_ CARRYB_11__3_ SUMB_11__3_ VDD VSS FA_X1 
XS2_11_2 ab_11__2_ CARRYB_10__2_ SUMB_10__3_ CARRYB_11__2_ SUMB_11__2_ VDD VSS FA_X1 
XS2_11_1 ab_11__1_ CARRYB_10__1_ SUMB_10__2_ CARRYB_11__1_ SUMB_11__1_ VDD VSS FA_X1 
XS1_11_0 ab_11__0_ CARRYB_10__0_ SUMB_10__1_ CARRYB_11__0_ A1_9_ VDD VSS FA_X1 
XS3_12_16 ab_12__16_ CARRYB_11__16_ ab_11__17_ CARRYB_12__16_ SUMB_12__16_ VDD VSS FA_X1 
XS2_12_15 ab_12__15_ CARRYB_11__15_ SUMB_11__16_ CARRYB_12__15_ SUMB_12__15_ VDD 
+ VSS FA_X1 
XS2_12_14 ab_12__14_ CARRYB_11__14_ SUMB_11__15_ CARRYB_12__14_ SUMB_12__14_ VDD 
+ VSS FA_X1 
XS2_12_13 ab_12__13_ CARRYB_11__13_ SUMB_11__14_ CARRYB_12__13_ SUMB_12__13_ VDD 
+ VSS FA_X1 
XS2_12_12 ab_12__12_ CARRYB_11__12_ SUMB_11__13_ CARRYB_12__12_ SUMB_12__12_ VDD 
+ VSS FA_X1 
XS2_12_11 ab_12__11_ CARRYB_11__11_ SUMB_11__12_ CARRYB_12__11_ SUMB_12__11_ VDD 
+ VSS FA_X1 
XS2_12_10 ab_12__10_ CARRYB_11__10_ SUMB_11__11_ CARRYB_12__10_ SUMB_12__10_ VDD 
+ VSS FA_X1 
XS2_12_9 ab_12__9_ CARRYB_11__9_ SUMB_11__10_ CARRYB_12__9_ SUMB_12__9_ VDD VSS FA_X1 
XS2_12_8 ab_12__8_ CARRYB_11__8_ SUMB_11__9_ CARRYB_12__8_ SUMB_12__8_ VDD VSS FA_X1 
XS2_12_7 ab_12__7_ CARRYB_11__7_ SUMB_11__8_ CARRYB_12__7_ SUMB_12__7_ VDD VSS FA_X1 
XS2_12_6 ab_12__6_ CARRYB_11__6_ SUMB_11__7_ CARRYB_12__6_ SUMB_12__6_ VDD VSS FA_X1 
XS2_12_5 ab_12__5_ CARRYB_11__5_ SUMB_11__6_ CARRYB_12__5_ SUMB_12__5_ VDD VSS FA_X1 
XS2_12_4 ab_12__4_ CARRYB_11__4_ SUMB_11__5_ CARRYB_12__4_ SUMB_12__4_ VDD VSS FA_X1 
XS2_12_3 ab_12__3_ CARRYB_11__3_ SUMB_11__4_ CARRYB_12__3_ SUMB_12__3_ VDD VSS FA_X1 
XS2_12_2 ab_12__2_ CARRYB_11__2_ SUMB_11__3_ CARRYB_12__2_ SUMB_12__2_ VDD VSS FA_X1 
XS2_12_1 ab_12__1_ CARRYB_11__1_ SUMB_11__2_ CARRYB_12__1_ SUMB_12__1_ VDD VSS FA_X1 
XS1_12_0 ab_12__0_ CARRYB_11__0_ SUMB_11__1_ CARRYB_12__0_ A1_10_ VDD VSS FA_X1 
XS3_13_16 ab_13__16_ CARRYB_12__16_ ab_12__17_ CARRYB_13__16_ SUMB_13__16_ VDD VSS FA_X1 
XS2_13_15 ab_13__15_ CARRYB_12__15_ SUMB_12__16_ CARRYB_13__15_ SUMB_13__15_ VDD 
+ VSS FA_X1 
XS2_13_14 ab_13__14_ CARRYB_12__14_ SUMB_12__15_ CARRYB_13__14_ SUMB_13__14_ VDD 
+ VSS FA_X1 
XS2_13_13 ab_13__13_ CARRYB_12__13_ SUMB_12__14_ CARRYB_13__13_ SUMB_13__13_ VDD 
+ VSS FA_X1 
XS2_13_12 ab_13__12_ CARRYB_12__12_ SUMB_12__13_ CARRYB_13__12_ SUMB_13__12_ VDD 
+ VSS FA_X1 
XS2_13_11 ab_13__11_ CARRYB_12__11_ SUMB_12__12_ CARRYB_13__11_ SUMB_13__11_ VDD 
+ VSS FA_X1 
XS2_13_10 ab_13__10_ CARRYB_12__10_ SUMB_12__11_ CARRYB_13__10_ SUMB_13__10_ VDD 
+ VSS FA_X1 
XS2_13_9 ab_13__9_ CARRYB_12__9_ SUMB_12__10_ CARRYB_13__9_ SUMB_13__9_ VDD VSS FA_X1 
XS2_13_8 ab_13__8_ CARRYB_12__8_ SUMB_12__9_ CARRYB_13__8_ SUMB_13__8_ VDD VSS FA_X1 
XS2_13_7 ab_13__7_ CARRYB_12__7_ SUMB_12__8_ CARRYB_13__7_ SUMB_13__7_ VDD VSS FA_X1 
XS2_13_6 ab_13__6_ CARRYB_12__6_ SUMB_12__7_ CARRYB_13__6_ SUMB_13__6_ VDD VSS FA_X1 
XS2_13_5 ab_13__5_ CARRYB_12__5_ SUMB_12__6_ CARRYB_13__5_ SUMB_13__5_ VDD VSS FA_X1 
XS2_13_4 ab_13__4_ CARRYB_12__4_ SUMB_12__5_ CARRYB_13__4_ SUMB_13__4_ VDD VSS FA_X1 
XS2_13_3 ab_13__3_ CARRYB_12__3_ SUMB_12__4_ CARRYB_13__3_ SUMB_13__3_ VDD VSS FA_X1 
XS2_13_2 ab_13__2_ CARRYB_12__2_ SUMB_12__3_ CARRYB_13__2_ SUMB_13__2_ VDD VSS FA_X1 
XS2_13_1 ab_13__1_ CARRYB_12__1_ SUMB_12__2_ CARRYB_13__1_ SUMB_13__1_ VDD VSS FA_X1 
XS1_13_0 ab_13__0_ CARRYB_12__0_ SUMB_12__1_ CARRYB_13__0_ A1_11_ VDD VSS FA_X1 
XS3_14_16 ab_14__16_ CARRYB_13__16_ ab_13__17_ CARRYB_14__16_ SUMB_14__16_ VDD VSS FA_X1 
XS2_14_15 ab_14__15_ CARRYB_13__15_ SUMB_13__16_ CARRYB_14__15_ SUMB_14__15_ VDD 
+ VSS FA_X1 
XS2_14_14 ab_14__14_ CARRYB_13__14_ SUMB_13__15_ CARRYB_14__14_ SUMB_14__14_ VDD 
+ VSS FA_X1 
XS2_14_13 ab_14__13_ CARRYB_13__13_ SUMB_13__14_ CARRYB_14__13_ SUMB_14__13_ VDD 
+ VSS FA_X1 
XS2_14_12 ab_14__12_ CARRYB_13__12_ SUMB_13__13_ CARRYB_14__12_ SUMB_14__12_ VDD 
+ VSS FA_X1 
XS2_14_11 ab_14__11_ CARRYB_13__11_ SUMB_13__12_ CARRYB_14__11_ SUMB_14__11_ VDD 
+ VSS FA_X1 
XS2_14_10 ab_14__10_ CARRYB_13__10_ SUMB_13__11_ CARRYB_14__10_ SUMB_14__10_ VDD 
+ VSS FA_X1 
XS2_14_9 ab_14__9_ CARRYB_13__9_ SUMB_13__10_ CARRYB_14__9_ SUMB_14__9_ VDD VSS FA_X1 
XS2_14_8 ab_14__8_ CARRYB_13__8_ SUMB_13__9_ CARRYB_14__8_ SUMB_14__8_ VDD VSS FA_X1 
XS2_14_7 ab_14__7_ CARRYB_13__7_ SUMB_13__8_ CARRYB_14__7_ SUMB_14__7_ VDD VSS FA_X1 
XS2_14_6 ab_14__6_ CARRYB_13__6_ SUMB_13__7_ CARRYB_14__6_ SUMB_14__6_ VDD VSS FA_X1 
XS2_14_5 ab_14__5_ CARRYB_13__5_ SUMB_13__6_ CARRYB_14__5_ SUMB_14__5_ VDD VSS FA_X1 
XS2_14_4 ab_14__4_ CARRYB_13__4_ SUMB_13__5_ CARRYB_14__4_ SUMB_14__4_ VDD VSS FA_X1 
XS2_14_3 ab_14__3_ CARRYB_13__3_ SUMB_13__4_ CARRYB_14__3_ SUMB_14__3_ VDD VSS FA_X1 
XS2_14_2 ab_14__2_ CARRYB_13__2_ SUMB_13__3_ CARRYB_14__2_ SUMB_14__2_ VDD VSS FA_X1 
XS2_14_1 ab_14__1_ CARRYB_13__1_ SUMB_13__2_ CARRYB_14__1_ SUMB_14__1_ VDD VSS FA_X1 
XS1_14_0 ab_14__0_ CARRYB_13__0_ SUMB_13__1_ CARRYB_14__0_ A1_12_ VDD VSS FA_X1 
XS14_17 n1 n85 ab_15__17_ CARRYB_15__17_ SUMB_15__17_ VDD VSS FA_X1 
XS5_16 ab_15__16_ CARRYB_14__16_ ab_14__17_ CARRYB_15__16_ SUMB_15__16_ VDD VSS FA_X1 
XS4_15 ab_15__15_ CARRYB_14__15_ SUMB_14__16_ CARRYB_15__15_ SUMB_15__15_ VDD VSS FA_X1 
XS4_14 ab_15__14_ CARRYB_14__14_ SUMB_14__15_ CARRYB_15__14_ SUMB_15__14_ VDD VSS FA_X1 
XS4_13 ab_15__13_ CARRYB_14__13_ SUMB_14__14_ CARRYB_15__13_ SUMB_15__13_ VDD VSS FA_X1 
XS4_12 ab_15__12_ CARRYB_14__12_ SUMB_14__13_ CARRYB_15__12_ SUMB_15__12_ VDD VSS FA_X1 
XS4_11 ab_15__11_ CARRYB_14__11_ SUMB_14__12_ CARRYB_15__11_ SUMB_15__11_ VDD VSS FA_X1 
XS4_10 ab_15__10_ CARRYB_14__10_ SUMB_14__11_ CARRYB_15__10_ SUMB_15__10_ VDD VSS FA_X1 
XS4_9 ab_15__9_ CARRYB_14__9_ SUMB_14__10_ CARRYB_15__9_ SUMB_15__9_ VDD VSS FA_X1 
XS4_8 ab_15__8_ CARRYB_14__8_ SUMB_14__9_ CARRYB_15__8_ SUMB_15__8_ VDD VSS FA_X1 
XS4_7 ab_15__7_ CARRYB_14__7_ SUMB_14__8_ CARRYB_15__7_ SUMB_15__7_ VDD VSS FA_X1 
XS4_6 ab_15__6_ CARRYB_14__6_ SUMB_14__7_ CARRYB_15__6_ SUMB_15__6_ VDD VSS FA_X1 
XS4_5 ab_15__5_ CARRYB_14__5_ SUMB_14__6_ CARRYB_15__5_ SUMB_15__5_ VDD VSS FA_X1 
XS4_4 ab_15__4_ CARRYB_14__4_ SUMB_14__5_ CARRYB_15__4_ SUMB_15__4_ VDD VSS FA_X1 
XS4_3 ab_15__3_ CARRYB_14__3_ SUMB_14__4_ CARRYB_15__3_ SUMB_15__3_ VDD VSS FA_X1 
XS4_2 ab_15__2_ CARRYB_14__2_ SUMB_14__3_ CARRYB_15__2_ SUMB_15__2_ VDD VSS FA_X1 
XS4_1 ab_15__1_ CARRYB_14__1_ SUMB_14__2_ CARRYB_15__1_ SUMB_15__1_ VDD VSS FA_X1 
XS4_0 ab_15__0_ CARRYB_14__0_ SUMB_14__1_ CARRYB_15__0_ SUMB_15__0_ VDD VSS FA_X1 
XS14_17_0 B[17] CARRYB_15__1_ SUMB_15__2_ A2_16_ A1_15_ VDD VSS FA_X1 
XS3_6_16 ab_6__16_ CARRYB_5__16_ ab_5__17_ CARRYB_6__16_ SUMB_6__16_ VDD VSS FA_X1 
XS2_6_15 ab_6__15_ CARRYB_5__15_ SUMB_5__16_ CARRYB_6__15_ SUMB_6__15_ VDD VSS FA_X1 
XS2_6_14 ab_6__14_ CARRYB_5__14_ SUMB_5__15_ CARRYB_6__14_ SUMB_6__14_ VDD VSS FA_X1 
XS2_6_13 ab_6__13_ CARRYB_5__13_ SUMB_5__14_ CARRYB_6__13_ SUMB_6__13_ VDD VSS FA_X1 
XS2_6_12 ab_6__12_ CARRYB_5__12_ SUMB_5__13_ CARRYB_6__12_ SUMB_6__12_ VDD VSS FA_X1 
XS2_6_11 ab_6__11_ CARRYB_5__11_ SUMB_5__12_ CARRYB_6__11_ SUMB_6__11_ VDD VSS FA_X1 
XS2_6_10 ab_6__10_ CARRYB_5__10_ SUMB_5__11_ CARRYB_6__10_ SUMB_6__10_ VDD VSS FA_X1 
XS2_6_9 ab_6__9_ CARRYB_5__9_ SUMB_5__10_ CARRYB_6__9_ SUMB_6__9_ VDD VSS FA_X1 
XS2_6_8 ab_6__8_ CARRYB_5__8_ SUMB_5__9_ CARRYB_6__8_ SUMB_6__8_ VDD VSS FA_X1 
XS2_6_7 ab_6__7_ CARRYB_5__7_ SUMB_5__8_ CARRYB_6__7_ SUMB_6__7_ VDD VSS FA_X1 
XS2_6_6 ab_6__6_ CARRYB_5__6_ SUMB_5__7_ CARRYB_6__6_ SUMB_6__6_ VDD VSS FA_X1 
XS2_6_5 ab_6__5_ CARRYB_5__5_ SUMB_5__6_ CARRYB_6__5_ SUMB_6__5_ VDD VSS FA_X1 
XS2_6_4 ab_6__4_ CARRYB_5__4_ SUMB_5__5_ CARRYB_6__4_ SUMB_6__4_ VDD VSS FA_X1 
XS2_6_3 ab_6__3_ CARRYB_5__3_ SUMB_5__4_ CARRYB_6__3_ SUMB_6__3_ VDD VSS FA_X1 
XS2_6_2 ab_6__2_ CARRYB_5__2_ SUMB_5__3_ CARRYB_6__2_ SUMB_6__2_ VDD VSS FA_X1 
XS2_6_1 ab_6__1_ CARRYB_5__1_ SUMB_5__2_ CARRYB_6__1_ SUMB_6__1_ VDD VSS FA_X1 
XS1_6_0 ab_6__0_ CARRYB_5__0_ SUMB_5__1_ CARRYB_6__0_ A1_4_ VDD VSS FA_X1 
XS3_7_16 ab_7__16_ CARRYB_6__16_ ab_6__17_ CARRYB_7__16_ SUMB_7__16_ VDD VSS FA_X1 
XS2_7_15 ab_7__15_ CARRYB_6__15_ SUMB_6__16_ CARRYB_7__15_ SUMB_7__15_ VDD VSS FA_X1 
XS2_7_14 ab_7__14_ CARRYB_6__14_ SUMB_6__15_ CARRYB_7__14_ SUMB_7__14_ VDD VSS FA_X1 
XS2_7_13 ab_7__13_ CARRYB_6__13_ SUMB_6__14_ CARRYB_7__13_ SUMB_7__13_ VDD VSS FA_X1 
XS2_7_12 ab_7__12_ CARRYB_6__12_ SUMB_6__13_ CARRYB_7__12_ SUMB_7__12_ VDD VSS FA_X1 
XS2_7_11 ab_7__11_ CARRYB_6__11_ SUMB_6__12_ CARRYB_7__11_ SUMB_7__11_ VDD VSS FA_X1 
XS2_7_10 ab_7__10_ CARRYB_6__10_ SUMB_6__11_ CARRYB_7__10_ SUMB_7__10_ VDD VSS FA_X1 
XS2_7_9 ab_7__9_ CARRYB_6__9_ SUMB_6__10_ CARRYB_7__9_ SUMB_7__9_ VDD VSS FA_X1 
XS2_7_8 ab_7__8_ CARRYB_6__8_ SUMB_6__9_ CARRYB_7__8_ SUMB_7__8_ VDD VSS FA_X1 
XS2_7_7 ab_7__7_ CARRYB_6__7_ SUMB_6__8_ CARRYB_7__7_ SUMB_7__7_ VDD VSS FA_X1 
XS2_7_6 ab_7__6_ CARRYB_6__6_ SUMB_6__7_ CARRYB_7__6_ SUMB_7__6_ VDD VSS FA_X1 
XS2_7_5 ab_7__5_ CARRYB_6__5_ SUMB_6__6_ CARRYB_7__5_ SUMB_7__5_ VDD VSS FA_X1 
XS2_7_4 ab_7__4_ CARRYB_6__4_ SUMB_6__5_ CARRYB_7__4_ SUMB_7__4_ VDD VSS FA_X1 
XS2_7_3 ab_7__3_ CARRYB_6__3_ SUMB_6__4_ CARRYB_7__3_ SUMB_7__3_ VDD VSS FA_X1 
XS2_7_2 ab_7__2_ CARRYB_6__2_ SUMB_6__3_ CARRYB_7__2_ SUMB_7__2_ VDD VSS FA_X1 
XS2_7_1 ab_7__1_ CARRYB_6__1_ SUMB_6__2_ CARRYB_7__1_ SUMB_7__1_ VDD VSS FA_X1 
XS1_7_0 ab_7__0_ CARRYB_6__0_ SUMB_6__1_ CARRYB_7__0_ A1_5_ VDD VSS FA_X1 
XS3_8_16 ab_8__16_ CARRYB_7__16_ ab_7__17_ CARRYB_8__16_ SUMB_8__16_ VDD VSS FA_X1 
XS2_8_15 ab_8__15_ CARRYB_7__15_ SUMB_7__16_ CARRYB_8__15_ SUMB_8__15_ VDD VSS FA_X1 
XS2_8_14 ab_8__14_ CARRYB_7__14_ SUMB_7__15_ CARRYB_8__14_ SUMB_8__14_ VDD VSS FA_X1 
XS2_8_13 ab_8__13_ CARRYB_7__13_ SUMB_7__14_ CARRYB_8__13_ SUMB_8__13_ VDD VSS FA_X1 
XS2_8_12 ab_8__12_ CARRYB_7__12_ SUMB_7__13_ CARRYB_8__12_ SUMB_8__12_ VDD VSS FA_X1 
XS2_8_11 ab_8__11_ CARRYB_7__11_ SUMB_7__12_ CARRYB_8__11_ SUMB_8__11_ VDD VSS FA_X1 
XS2_8_10 ab_8__10_ CARRYB_7__10_ SUMB_7__11_ CARRYB_8__10_ SUMB_8__10_ VDD VSS FA_X1 
XS2_8_9 ab_8__9_ CARRYB_7__9_ SUMB_7__10_ CARRYB_8__9_ SUMB_8__9_ VDD VSS FA_X1 
XS2_8_8 ab_8__8_ CARRYB_7__8_ SUMB_7__9_ CARRYB_8__8_ SUMB_8__8_ VDD VSS FA_X1 
XS2_8_7 ab_8__7_ CARRYB_7__7_ SUMB_7__8_ CARRYB_8__7_ SUMB_8__7_ VDD VSS FA_X1 
XS2_8_6 ab_8__6_ CARRYB_7__6_ SUMB_7__7_ CARRYB_8__6_ SUMB_8__6_ VDD VSS FA_X1 
XS2_8_5 ab_8__5_ CARRYB_7__5_ SUMB_7__6_ CARRYB_8__5_ SUMB_8__5_ VDD VSS FA_X1 
XS2_8_4 ab_8__4_ CARRYB_7__4_ SUMB_7__5_ CARRYB_8__4_ SUMB_8__4_ VDD VSS FA_X1 
XS2_8_3 ab_8__3_ CARRYB_7__3_ SUMB_7__4_ CARRYB_8__3_ SUMB_8__3_ VDD VSS FA_X1 
XS2_8_2 ab_8__2_ CARRYB_7__2_ SUMB_7__3_ CARRYB_8__2_ SUMB_8__2_ VDD VSS FA_X1 
XS2_8_1 ab_8__1_ CARRYB_7__1_ SUMB_7__2_ CARRYB_8__1_ SUMB_8__1_ VDD VSS FA_X1 
XS1_8_0 ab_8__0_ CARRYB_7__0_ SUMB_7__1_ CARRYB_8__0_ A1_6_ VDD VSS FA_X1 
XS3_9_16 ab_9__16_ CARRYB_8__16_ ab_8__17_ CARRYB_9__16_ SUMB_9__16_ VDD VSS FA_X1 
XS2_9_15 ab_9__15_ CARRYB_8__15_ SUMB_8__16_ CARRYB_9__15_ SUMB_9__15_ VDD VSS FA_X1 
XS2_9_14 ab_9__14_ CARRYB_8__14_ SUMB_8__15_ CARRYB_9__14_ SUMB_9__14_ VDD VSS FA_X1 
XS2_9_13 ab_9__13_ CARRYB_8__13_ SUMB_8__14_ CARRYB_9__13_ SUMB_9__13_ VDD VSS FA_X1 
XS2_9_12 ab_9__12_ CARRYB_8__12_ SUMB_8__13_ CARRYB_9__12_ SUMB_9__12_ VDD VSS FA_X1 
XS2_9_11 ab_9__11_ CARRYB_8__11_ SUMB_8__12_ CARRYB_9__11_ SUMB_9__11_ VDD VSS FA_X1 
XS2_9_10 ab_9__10_ CARRYB_8__10_ SUMB_8__11_ CARRYB_9__10_ SUMB_9__10_ VDD VSS FA_X1 
XS2_9_9 ab_9__9_ CARRYB_8__9_ SUMB_8__10_ CARRYB_9__9_ SUMB_9__9_ VDD VSS FA_X1 
XS2_9_8 ab_9__8_ CARRYB_8__8_ SUMB_8__9_ CARRYB_9__8_ SUMB_9__8_ VDD VSS FA_X1 
XS2_9_7 ab_9__7_ CARRYB_8__7_ SUMB_8__8_ CARRYB_9__7_ SUMB_9__7_ VDD VSS FA_X1 
XS2_9_6 ab_9__6_ CARRYB_8__6_ SUMB_8__7_ CARRYB_9__6_ SUMB_9__6_ VDD VSS FA_X1 
XS2_9_5 ab_9__5_ CARRYB_8__5_ SUMB_8__6_ CARRYB_9__5_ SUMB_9__5_ VDD VSS FA_X1 
XS2_9_4 ab_9__4_ CARRYB_8__4_ SUMB_8__5_ CARRYB_9__4_ SUMB_9__4_ VDD VSS FA_X1 
XS2_9_3 ab_9__3_ CARRYB_8__3_ SUMB_8__4_ CARRYB_9__3_ SUMB_9__3_ VDD VSS FA_X1 
XS2_9_2 ab_9__2_ CARRYB_8__2_ SUMB_8__3_ CARRYB_9__2_ SUMB_9__2_ VDD VSS FA_X1 
XS2_9_1 ab_9__1_ CARRYB_8__1_ SUMB_8__2_ CARRYB_9__1_ SUMB_9__1_ VDD VSS FA_X1 
XS1_9_0 ab_9__0_ CARRYB_8__0_ SUMB_8__1_ CARRYB_9__0_ A1_7_ VDD VSS FA_X1 
XS3_10_16 ab_10__16_ CARRYB_9__16_ ab_9__17_ CARRYB_10__16_ SUMB_10__16_ VDD VSS FA_X1 
XS2_10_15 ab_10__15_ CARRYB_9__15_ SUMB_9__16_ CARRYB_10__15_ SUMB_10__15_ VDD VSS FA_X1 
XS2_10_14 ab_10__14_ CARRYB_9__14_ SUMB_9__15_ CARRYB_10__14_ SUMB_10__14_ VDD VSS FA_X1 
XS2_10_13 ab_10__13_ CARRYB_9__13_ SUMB_9__14_ CARRYB_10__13_ SUMB_10__13_ VDD VSS FA_X1 
XS2_10_12 ab_10__12_ CARRYB_9__12_ SUMB_9__13_ CARRYB_10__12_ SUMB_10__12_ VDD VSS FA_X1 
XS2_10_11 ab_10__11_ CARRYB_9__11_ SUMB_9__12_ CARRYB_10__11_ SUMB_10__11_ VDD VSS FA_X1 
XS2_10_10 ab_10__10_ CARRYB_9__10_ SUMB_9__11_ CARRYB_10__10_ SUMB_10__10_ VDD VSS FA_X1 
XS2_10_9 ab_10__9_ CARRYB_9__9_ SUMB_9__10_ CARRYB_10__9_ SUMB_10__9_ VDD VSS FA_X1 
XS2_10_8 ab_10__8_ CARRYB_9__8_ SUMB_9__9_ CARRYB_10__8_ SUMB_10__8_ VDD VSS FA_X1 
XS2_10_7 ab_10__7_ CARRYB_9__7_ SUMB_9__8_ CARRYB_10__7_ SUMB_10__7_ VDD VSS FA_X1 
XS2_10_6 ab_10__6_ CARRYB_9__6_ SUMB_9__7_ CARRYB_10__6_ SUMB_10__6_ VDD VSS FA_X1 
XS2_10_5 ab_10__5_ CARRYB_9__5_ SUMB_9__6_ CARRYB_10__5_ SUMB_10__5_ VDD VSS FA_X1 
XS2_10_4 ab_10__4_ CARRYB_9__4_ SUMB_9__5_ CARRYB_10__4_ SUMB_10__4_ VDD VSS FA_X1 
XS2_10_3 ab_10__3_ CARRYB_9__3_ SUMB_9__4_ CARRYB_10__3_ SUMB_10__3_ VDD VSS FA_X1 
XS2_10_2 ab_10__2_ CARRYB_9__2_ SUMB_9__3_ CARRYB_10__2_ SUMB_10__2_ VDD VSS FA_X1 
XS2_10_1 ab_10__1_ CARRYB_9__1_ SUMB_9__2_ CARRYB_10__1_ SUMB_10__1_ VDD VSS FA_X1 
XS1_10_0 ab_10__0_ CARRYB_9__0_ SUMB_9__1_ CARRYB_10__0_ A1_8_ VDD VSS FA_X1 
XS3_11_16 ab_11__16_ CARRYB_10__16_ ab_10__17_ CARRYB_11__16_ SUMB_11__16_ VDD VSS FA_X1 
XS2_11_15 ab_11__15_ CARRYB_10__15_ SUMB_10__16_ CARRYB_11__15_ SUMB_11__15_ VDD 
+ VSS FA_X1 
XS2_11_14 ab_11__14_ CARRYB_10__14_ SUMB_10__15_ CARRYB_11__14_ SUMB_11__14_ VDD 
+ VSS FA_X1 
XS2_11_13 ab_11__13_ CARRYB_10__13_ SUMB_10__14_ CARRYB_11__13_ SUMB_11__13_ VDD 
+ VSS FA_X1 
XS2_11_12 ab_11__12_ CARRYB_10__12_ SUMB_10__13_ CARRYB_11__12_ SUMB_11__12_ VDD 
+ VSS FA_X1 
XS2_11_11 ab_11__11_ CARRYB_10__11_ SUMB_10__12_ CARRYB_11__11_ SUMB_11__11_ VDD 
+ VSS FA_X1 
XS2_11_10 ab_11__10_ CARRYB_10__10_ SUMB_10__11_ CARRYB_11__10_ SUMB_11__10_ VDD 
+ VSS FA_X1 
XS2_11_9 ab_11__9_ CARRYB_10__9_ SUMB_10__10_ CARRYB_11__9_ SUMB_11__9_ VDD VSS FA_X1 
XU26 ab_1__8_ ab_0__9_ n26 VDD VSS XOR2_X1 
XU25 ab_1__9_ ab_0__10_ n25 VDD VSS XOR2_X1 
XU24 ab_1__10_ ab_0__11_ n24 VDD VSS XOR2_X1 
XU23 ab_1__11_ ab_0__12_ n23 VDD VSS XOR2_X1 
XU22 ab_1__12_ ab_0__13_ n22 VDD VSS XOR2_X1 
XU21 ab_1__13_ ab_0__14_ n21 VDD VSS XOR2_X1 
XU20 ab_1__14_ ab_0__15_ n20 VDD VSS XOR2_X1 
XU19 ab_1__15_ ab_0__16_ n19 VDD VSS XOR2_X1 
XU18 ab_0__17_ ab_1__16_ n18 VDD VSS AND2_X1 
XU17 ab_0__1_ ab_1__0_ n17 VDD VSS AND2_X1 
XU16 ab_0__2_ ab_1__1_ n16 VDD VSS AND2_X1 
XU15 ab_0__3_ ab_1__2_ n15 VDD VSS AND2_X1 
XU14 ab_0__4_ ab_1__3_ n14 VDD VSS AND2_X1 
XU13 ab_0__5_ ab_1__4_ n13 VDD VSS AND2_X1 
XU12 ab_0__6_ ab_1__5_ n12 VDD VSS AND2_X1 
XU11 ab_0__7_ ab_1__6_ n11 VDD VSS AND2_X1 
XU10 ab_0__8_ ab_1__7_ n10 VDD VSS AND2_X1 
XU9 ab_0__9_ ab_1__8_ n9 VDD VSS AND2_X1 
XU8 ab_0__10_ ab_1__9_ n8 VDD VSS AND2_X1 
XU7 ab_0__11_ ab_1__10_ n7 VDD VSS AND2_X1 
XU6 ab_0__12_ ab_1__11_ n6 VDD VSS AND2_X1 
XU5 ab_0__13_ ab_1__12_ n5 VDD VSS AND2_X1 
XU4 ab_0__14_ ab_1__13_ n4 VDD VSS AND2_X1 
XU3 ab_0__15_ ab_1__14_ n3 VDD VSS AND2_X1 
XU2 ab_0__16_ ab_1__15_ n2 VDD VSS AND2_X1 
XS3_2_16 ab_2__16_ n18 ab_1__17_ CARRYB_2__16_ SUMB_2__16_ VDD VSS FA_X1 
XS2_2_15 ab_2__15_ n2 n32 CARRYB_2__15_ SUMB_2__15_ VDD VSS FA_X1 
XS2_2_14 ab_2__14_ n3 n19 CARRYB_2__14_ SUMB_2__14_ VDD VSS FA_X1 
XS2_2_13 ab_2__13_ n4 n20 CARRYB_2__13_ SUMB_2__13_ VDD VSS FA_X1 
XS2_2_12 ab_2__12_ n5 n21 CARRYB_2__12_ SUMB_2__12_ VDD VSS FA_X1 
XS2_2_11 ab_2__11_ n6 n22 CARRYB_2__11_ SUMB_2__11_ VDD VSS FA_X1 
XS2_2_10 ab_2__10_ n7 n23 CARRYB_2__10_ SUMB_2__10_ VDD VSS FA_X1 
XS2_2_9 ab_2__9_ n8 n24 CARRYB_2__9_ SUMB_2__9_ VDD VSS FA_X1 
XS2_2_8 ab_2__8_ n9 n25 CARRYB_2__8_ SUMB_2__8_ VDD VSS FA_X1 
XS2_2_7 ab_2__7_ n10 n26 CARRYB_2__7_ SUMB_2__7_ VDD VSS FA_X1 
XS2_2_6 ab_2__6_ n11 n27 CARRYB_2__6_ SUMB_2__6_ VDD VSS FA_X1 
XS2_2_5 ab_2__5_ n12 n28 CARRYB_2__5_ SUMB_2__5_ VDD VSS FA_X1 
XS2_2_4 ab_2__4_ n13 n29 CARRYB_2__4_ SUMB_2__4_ VDD VSS FA_X1 
XS2_2_3 ab_2__3_ n14 n30 CARRYB_2__3_ SUMB_2__3_ VDD VSS FA_X1 
XS2_2_2 ab_2__2_ n15 n31 CARRYB_2__2_ SUMB_2__2_ VDD VSS FA_X1 
XS2_2_1 ab_2__1_ n16 n33 CARRYB_2__1_ SUMB_2__1_ VDD VSS FA_X1 
XS1_2_0 ab_2__0_ n17 n34 CARRYB_2__0_ A1_0_ VDD VSS FA_X1 
XS3_3_16 ab_3__16_ CARRYB_2__16_ ab_2__17_ CARRYB_3__16_ SUMB_3__16_ VDD VSS FA_X1 
XS2_3_15 ab_3__15_ CARRYB_2__15_ SUMB_2__16_ CARRYB_3__15_ SUMB_3__15_ VDD VSS FA_X1 
XS2_3_14 ab_3__14_ CARRYB_2__14_ SUMB_2__15_ CARRYB_3__14_ SUMB_3__14_ VDD VSS FA_X1 
XS2_3_13 ab_3__13_ CARRYB_2__13_ SUMB_2__14_ CARRYB_3__13_ SUMB_3__13_ VDD VSS FA_X1 
XS2_3_12 ab_3__12_ CARRYB_2__12_ SUMB_2__13_ CARRYB_3__12_ SUMB_3__12_ VDD VSS FA_X1 
XS2_3_11 ab_3__11_ CARRYB_2__11_ SUMB_2__12_ CARRYB_3__11_ SUMB_3__11_ VDD VSS FA_X1 
XS2_3_10 ab_3__10_ CARRYB_2__10_ SUMB_2__11_ CARRYB_3__10_ SUMB_3__10_ VDD VSS FA_X1 
XS2_3_9 ab_3__9_ CARRYB_2__9_ SUMB_2__10_ CARRYB_3__9_ SUMB_3__9_ VDD VSS FA_X1 
XS2_3_8 ab_3__8_ CARRYB_2__8_ SUMB_2__9_ CARRYB_3__8_ SUMB_3__8_ VDD VSS FA_X1 
XS2_3_7 ab_3__7_ CARRYB_2__7_ SUMB_2__8_ CARRYB_3__7_ SUMB_3__7_ VDD VSS FA_X1 
XS2_3_6 ab_3__6_ CARRYB_2__6_ SUMB_2__7_ CARRYB_3__6_ SUMB_3__6_ VDD VSS FA_X1 
XS2_3_5 ab_3__5_ CARRYB_2__5_ SUMB_2__6_ CARRYB_3__5_ SUMB_3__5_ VDD VSS FA_X1 
XS2_3_4 ab_3__4_ CARRYB_2__4_ SUMB_2__5_ CARRYB_3__4_ SUMB_3__4_ VDD VSS FA_X1 
XS2_3_3 ab_3__3_ CARRYB_2__3_ SUMB_2__4_ CARRYB_3__3_ SUMB_3__3_ VDD VSS FA_X1 
XS2_3_2 ab_3__2_ CARRYB_2__2_ SUMB_2__3_ CARRYB_3__2_ SUMB_3__2_ VDD VSS FA_X1 
XS2_3_1 ab_3__1_ CARRYB_2__1_ SUMB_2__2_ CARRYB_3__1_ SUMB_3__1_ VDD VSS FA_X1 
XS1_3_0 ab_3__0_ CARRYB_2__0_ SUMB_2__1_ CARRYB_3__0_ A1_1_ VDD VSS FA_X1 
XS3_4_16 ab_4__16_ CARRYB_3__16_ ab_3__17_ CARRYB_4__16_ SUMB_4__16_ VDD VSS FA_X1 
XS2_4_15 ab_4__15_ CARRYB_3__15_ SUMB_3__16_ CARRYB_4__15_ SUMB_4__15_ VDD VSS FA_X1 
XS2_4_14 ab_4__14_ CARRYB_3__14_ SUMB_3__15_ CARRYB_4__14_ SUMB_4__14_ VDD VSS FA_X1 
XS2_4_13 ab_4__13_ CARRYB_3__13_ SUMB_3__14_ CARRYB_4__13_ SUMB_4__13_ VDD VSS FA_X1 
XS2_4_12 ab_4__12_ CARRYB_3__12_ SUMB_3__13_ CARRYB_4__12_ SUMB_4__12_ VDD VSS FA_X1 
XS2_4_11 ab_4__11_ CARRYB_3__11_ SUMB_3__12_ CARRYB_4__11_ SUMB_4__11_ VDD VSS FA_X1 
XS2_4_10 ab_4__10_ CARRYB_3__10_ SUMB_3__11_ CARRYB_4__10_ SUMB_4__10_ VDD VSS FA_X1 
XS2_4_9 ab_4__9_ CARRYB_3__9_ SUMB_3__10_ CARRYB_4__9_ SUMB_4__9_ VDD VSS FA_X1 
XS2_4_8 ab_4__8_ CARRYB_3__8_ SUMB_3__9_ CARRYB_4__8_ SUMB_4__8_ VDD VSS FA_X1 
XS2_4_7 ab_4__7_ CARRYB_3__7_ SUMB_3__8_ CARRYB_4__7_ SUMB_4__7_ VDD VSS FA_X1 
XS2_4_6 ab_4__6_ CARRYB_3__6_ SUMB_3__7_ CARRYB_4__6_ SUMB_4__6_ VDD VSS FA_X1 
XS2_4_5 ab_4__5_ CARRYB_3__5_ SUMB_3__6_ CARRYB_4__5_ SUMB_4__5_ VDD VSS FA_X1 
XS2_4_4 ab_4__4_ CARRYB_3__4_ SUMB_3__5_ CARRYB_4__4_ SUMB_4__4_ VDD VSS FA_X1 
XS2_4_3 ab_4__3_ CARRYB_3__3_ SUMB_3__4_ CARRYB_4__3_ SUMB_4__3_ VDD VSS FA_X1 
XS2_4_2 ab_4__2_ CARRYB_3__2_ SUMB_3__3_ CARRYB_4__2_ SUMB_4__2_ VDD VSS FA_X1 
XS2_4_1 ab_4__1_ CARRYB_3__1_ SUMB_3__2_ CARRYB_4__1_ SUMB_4__1_ VDD VSS FA_X1 
XS1_4_0 ab_4__0_ CARRYB_3__0_ SUMB_3__1_ CARRYB_4__0_ A1_2_ VDD VSS FA_X1 
XS3_5_16 ab_5__16_ CARRYB_4__16_ ab_4__17_ CARRYB_5__16_ SUMB_5__16_ VDD VSS FA_X1 
XS2_5_15 ab_5__15_ CARRYB_4__15_ SUMB_4__16_ CARRYB_5__15_ SUMB_5__15_ VDD VSS FA_X1 
XS2_5_14 ab_5__14_ CARRYB_4__14_ SUMB_4__15_ CARRYB_5__14_ SUMB_5__14_ VDD VSS FA_X1 
XS2_5_13 ab_5__13_ CARRYB_4__13_ SUMB_4__14_ CARRYB_5__13_ SUMB_5__13_ VDD VSS FA_X1 
XS2_5_12 ab_5__12_ CARRYB_4__12_ SUMB_4__13_ CARRYB_5__12_ SUMB_5__12_ VDD VSS FA_X1 
XS2_5_11 ab_5__11_ CARRYB_4__11_ SUMB_4__12_ CARRYB_5__11_ SUMB_5__11_ VDD VSS FA_X1 
XS2_5_10 ab_5__10_ CARRYB_4__10_ SUMB_4__11_ CARRYB_5__10_ SUMB_5__10_ VDD VSS FA_X1 
XS2_5_9 ab_5__9_ CARRYB_4__9_ SUMB_4__10_ CARRYB_5__9_ SUMB_5__9_ VDD VSS FA_X1 
XS2_5_8 ab_5__8_ CARRYB_4__8_ SUMB_4__9_ CARRYB_5__8_ SUMB_5__8_ VDD VSS FA_X1 
XS2_5_7 ab_5__7_ CARRYB_4__7_ SUMB_4__8_ CARRYB_5__7_ SUMB_5__7_ VDD VSS FA_X1 
XS2_5_6 ab_5__6_ CARRYB_4__6_ SUMB_4__7_ CARRYB_5__6_ SUMB_5__6_ VDD VSS FA_X1 
XS2_5_5 ab_5__5_ CARRYB_4__5_ SUMB_4__6_ CARRYB_5__5_ SUMB_5__5_ VDD VSS FA_X1 
XS2_5_4 ab_5__4_ CARRYB_4__4_ SUMB_4__5_ CARRYB_5__4_ SUMB_5__4_ VDD VSS FA_X1 
XS2_5_3 ab_5__3_ CARRYB_4__3_ SUMB_4__4_ CARRYB_5__3_ SUMB_5__3_ VDD VSS FA_X1 
XS2_5_2 ab_5__2_ CARRYB_4__2_ SUMB_4__3_ CARRYB_5__2_ SUMB_5__2_ VDD VSS FA_X1 
XS2_5_1 ab_5__1_ CARRYB_4__1_ SUMB_4__2_ CARRYB_5__1_ SUMB_5__1_ VDD VSS FA_X1 
XS1_5_0 ab_5__0_ CARRYB_4__0_ SUMB_4__1_ CARRYB_5__0_ A1_3_ VDD VSS FA_X1 
XU119 n75 n90 ab_9__12_ VDD VSS NOR2_X1 
XU118 n75 n89 ab_9__13_ VDD VSS NOR2_X1 
XU117 n75 n88 ab_9__14_ VDD VSS NOR2_X1 
XU116 n75 n87 ab_9__15_ VDD VSS NOR2_X1 
XU115 n75 n86 ab_9__16_ VDD VSS NOR2_X1 
XU114 A[9] n85 ab_9__17_ VDD VSS NOR2_X1 
XU113 n75 n101 ab_9__1_ VDD VSS NOR2_X1 
XU112 n75 n100 ab_9__2_ VDD VSS NOR2_X1 
XU111 n75 n99 ab_9__3_ VDD VSS NOR2_X1 
XU110 n75 n98 ab_9__4_ VDD VSS NOR2_X1 
XU109 n75 n97 ab_9__5_ VDD VSS NOR2_X1 
XU108 n75 n96 ab_9__6_ VDD VSS NOR2_X1 
XU107 n75 n95 ab_9__7_ VDD VSS NOR2_X1 
XU106 n75 n94 ab_9__8_ VDD VSS NOR2_X1 
XU105 n75 n93 ab_9__9_ VDD VSS NOR2_X1 
XU103 B[0] n102 VDD VSS INV_X1 
XU102 B[1] n101 VDD VSS INV_X1 
XU101 A[15] SUMB_15__0_ n69 VDD VSS XOR2_X1 
XU100 B[2] n100 VDD VSS INV_X1 
XU99 B[3] n99 VDD VSS INV_X1 
XU98 B[4] n98 VDD VSS INV_X1 
XU97 B[5] n97 VDD VSS INV_X1 
XU96 B[6] n96 VDD VSS INV_X1 
XU95 B[7] n95 VDD VSS INV_X1 
XU94 B[8] n94 VDD VSS INV_X1 
XU93 B[9] n93 VDD VSS INV_X1 
XU92 B[10] n92 VDD VSS INV_X1 
XU91 B[11] n91 VDD VSS INV_X1 
XU90 B[12] n90 VDD VSS INV_X1 
XU89 A[15] SUMB_15__0_ n68 VDD VSS AND2_X1 
XU88 B[13] n89 VDD VSS INV_X1 
XU87 B[14] n88 VDD VSS INV_X1 
XU86 B[15] n87 VDD VSS INV_X1 
XU85 B[16] n86 VDD VSS INV_X1 
XU84 B[17] n85 VDD VSS INV_X1 
XU83 A[0] n84 VDD VSS INV_X1 
XU82 A[1] n83 VDD VSS INV_X1 
XU81 A[2] n82 VDD VSS INV_X1 
XU80 A[3] n81 VDD VSS INV_X1 
XU79 A[4] n80 VDD VSS INV_X1 
XU78 A[5] n79 VDD VSS INV_X1 
XU77 A[6] n78 VDD VSS INV_X1 
XU76 A[7] n77 VDD VSS INV_X1 
XU75 A[8] n76 VDD VSS INV_X1 
XU74 A[9] n75 VDD VSS INV_X1 
XU73 A[10] n74 VDD VSS INV_X1 
XU72 A[11] n73 VDD VSS INV_X1 
XU71 A[12] n72 VDD VSS INV_X1 
XU70 A[13] n71 VDD VSS INV_X1 
XU69 A[14] n35 VDD VSS INV_X1 
XU68 CARRYB_15__15_ SUMB_15__16_ n67 VDD VSS XOR2_X1 
XU67 CARRYB_15__13_ SUMB_15__14_ n66 VDD VSS XOR2_X1 
XU66 CARRYB_15__11_ SUMB_15__12_ n65 VDD VSS XOR2_X1 
XU65 CARRYB_15__9_ SUMB_15__10_ n64 VDD VSS XOR2_X1 
XU64 CARRYB_15__7_ SUMB_15__8_ n63 VDD VSS XOR2_X1 
XU63 CARRYB_15__5_ SUMB_15__6_ n62 VDD VSS XOR2_X1 
XU62 CARRYB_15__15_ SUMB_15__16_ n61 VDD VSS AND2_X1 
XU61 CARRYB_15__14_ SUMB_15__15_ n60 VDD VSS AND2_X1 
XU60 CARRYB_15__13_ SUMB_15__14_ n59 VDD VSS AND2_X1 
XU59 CARRYB_15__12_ SUMB_15__13_ n58 VDD VSS AND2_X1 
XU58 CARRYB_15__11_ SUMB_15__12_ n57 VDD VSS AND2_X1 
XU57 CARRYB_15__10_ SUMB_15__11_ n56 VDD VSS AND2_X1 
XU56 CARRYB_15__9_ SUMB_15__10_ n55 VDD VSS AND2_X1 
XU55 CARRYB_15__8_ SUMB_15__9_ n54 VDD VSS AND2_X1 
XU54 CARRYB_15__7_ SUMB_15__8_ n53 VDD VSS AND2_X1 
XU53 CARRYB_15__6_ SUMB_15__7_ n52 VDD VSS AND2_X1 
XU52 CARRYB_15__5_ SUMB_15__6_ n51 VDD VSS AND2_X1 
XU51 CARRYB_15__4_ SUMB_15__5_ n50 VDD VSS AND2_X1 
XU50 CARRYB_15__16_ SUMB_15__17_ n49 VDD VSS AND2_X1 
XU49 CARRYB_15__16_ SUMB_15__17_ n48 VDD VSS XOR2_X1 
XU48 CARRYB_15__14_ SUMB_15__15_ n47 VDD VSS XOR2_X1 
XU47 CARRYB_15__12_ SUMB_15__13_ n46 VDD VSS XOR2_X1 
XU46 CARRYB_15__10_ SUMB_15__11_ n45 VDD VSS XOR2_X1 
XU45 CARRYB_15__8_ SUMB_15__9_ n44 VDD VSS XOR2_X1 
XU44 CARRYB_15__6_ SUMB_15__7_ n43 VDD VSS XOR2_X1 
XU43 CARRYB_15__3_ SUMB_15__4_ n42 VDD VSS XOR2_X1 
XU42 CARRYB_15__3_ SUMB_15__4_ n41 VDD VSS AND2_X1 
XU41 CARRYB_15__2_ SUMB_15__3_ n40 VDD VSS AND2_X1 
XU40 CARRYB_15__0_ SUMB_15__1_ n39 VDD VSS AND2_X1 
XU39 CARRYB_15__0_ SUMB_15__1_ n38 VDD VSS XOR2_X1 
XU38 CARRYB_15__4_ SUMB_15__5_ n37 VDD VSS XOR2_X1 
XU37 CARRYB_15__2_ SUMB_15__3_ n36 VDD VSS XOR2_X1 
XU36 ab_1__0_ ab_0__1_ n158 VDD VSS XOR2_X1 
XU35 CARRYB_15__17_ n70 VDD VSS INV_X1 
XU34 ab_1__1_ ab_0__2_ n34 VDD VSS XOR2_X1 
XU33 ab_1__2_ ab_0__3_ n33 VDD VSS XOR2_X1 
XU32 ab_1__16_ ab_0__17_ n32 VDD VSS XOR2_X1 
XU31 ab_1__3_ ab_0__4_ n31 VDD VSS XOR2_X1 
XU30 ab_1__4_ ab_0__5_ n30 VDD VSS XOR2_X1 
XU29 ab_1__5_ ab_0__6_ n29 VDD VSS XOR2_X1 
XU28 ab_1__6_ ab_0__7_ n28 VDD VSS XOR2_X1 
XU27 ab_1__7_ ab_0__8_ n27 VDD VSS XOR2_X1 
XU212 n156 n80 ab_4__0_ VDD VSS NOR2_X1 
XU211 n92 n80 ab_4__10_ VDD VSS NOR2_X1 
XU210 n91 n80 ab_4__11_ VDD VSS NOR2_X1 
XU209 n90 n80 ab_4__12_ VDD VSS NOR2_X1 
XU208 n89 n80 ab_4__13_ VDD VSS NOR2_X1 
XU207 n88 n80 ab_4__14_ VDD VSS NOR2_X1 
XU206 n87 n80 ab_4__15_ VDD VSS NOR2_X1 
XU205 n86 n80 ab_4__16_ VDD VSS NOR2_X1 
XU204 A[4] n85 ab_4__17_ VDD VSS NOR2_X1 
XU203 n101 n80 ab_4__1_ VDD VSS NOR2_X1 
XU202 n100 n80 ab_4__2_ VDD VSS NOR2_X1 
XU201 n99 n80 ab_4__3_ VDD VSS NOR2_X1 
XU200 n98 n80 ab_4__4_ VDD VSS NOR2_X1 
XU199 n97 n80 ab_4__5_ VDD VSS NOR2_X1 
XU198 n96 n80 ab_4__6_ VDD VSS NOR2_X1 
XU197 n95 n80 ab_4__7_ VDD VSS NOR2_X1 
XU196 n94 n80 ab_4__8_ VDD VSS NOR2_X1 
XU195 n93 n80 ab_4__9_ VDD VSS NOR2_X1 
XU194 n156 n79 ab_5__0_ VDD VSS NOR2_X1 
XU193 n92 n79 ab_5__10_ VDD VSS NOR2_X1 
XU192 n91 n79 ab_5__11_ VDD VSS NOR2_X1 
XU191 n90 n79 ab_5__12_ VDD VSS NOR2_X1 
XU190 n89 n79 ab_5__13_ VDD VSS NOR2_X1 
XU189 n88 n79 ab_5__14_ VDD VSS NOR2_X1 
XU188 n87 n79 ab_5__15_ VDD VSS NOR2_X1 
XU187 n86 n79 ab_5__16_ VDD VSS NOR2_X1 
XU186 A[5] n85 ab_5__17_ VDD VSS NOR2_X1 
XU185 n101 n79 ab_5__1_ VDD VSS NOR2_X1 
XU184 n100 n79 ab_5__2_ VDD VSS NOR2_X1 
XU183 n99 n79 ab_5__3_ VDD VSS NOR2_X1 
XU182 n98 n79 ab_5__4_ VDD VSS NOR2_X1 
XU181 n97 n79 ab_5__5_ VDD VSS NOR2_X1 
XU180 n96 n79 ab_5__6_ VDD VSS NOR2_X1 
XU179 n95 n79 ab_5__7_ VDD VSS NOR2_X1 
XU178 n94 n79 ab_5__8_ VDD VSS NOR2_X1 
XU177 n93 n79 ab_5__9_ VDD VSS NOR2_X1 
XU176 n156 n78 ab_6__0_ VDD VSS NOR2_X1 
XU175 n92 n78 ab_6__10_ VDD VSS NOR2_X1 
XU174 n91 n78 ab_6__11_ VDD VSS NOR2_X1 
XU173 n90 n78 ab_6__12_ VDD VSS NOR2_X1 
XU172 n89 n78 ab_6__13_ VDD VSS NOR2_X1 
XU171 n88 n78 ab_6__14_ VDD VSS NOR2_X1 
XU170 n87 n78 ab_6__15_ VDD VSS NOR2_X1 
XU169 n86 n78 ab_6__16_ VDD VSS NOR2_X1 
XU168 A[6] n85 ab_6__17_ VDD VSS NOR2_X1 
XU167 n101 n78 ab_6__1_ VDD VSS NOR2_X1 
XU166 n100 n78 ab_6__2_ VDD VSS NOR2_X1 
XU165 n99 n78 ab_6__3_ VDD VSS NOR2_X1 
XU164 n98 n78 ab_6__4_ VDD VSS NOR2_X1 
XU163 n97 n78 ab_6__5_ VDD VSS NOR2_X1 
XU162 n96 n78 ab_6__6_ VDD VSS NOR2_X1 
XU161 n95 n78 ab_6__7_ VDD VSS NOR2_X1 
XU160 n94 n78 ab_6__8_ VDD VSS NOR2_X1 
XU159 n93 n78 ab_6__9_ VDD VSS NOR2_X1 
XU158 n156 n77 ab_7__0_ VDD VSS NOR2_X1 
XU157 n92 n77 ab_7__10_ VDD VSS NOR2_X1 
XU156 n91 n77 ab_7__11_ VDD VSS NOR2_X1 
XU155 n90 n77 ab_7__12_ VDD VSS NOR2_X1 
XU154 n89 n77 ab_7__13_ VDD VSS NOR2_X1 
XU153 n88 n77 ab_7__14_ VDD VSS NOR2_X1 
XU152 n87 n77 ab_7__15_ VDD VSS NOR2_X1 
XU151 n86 n77 ab_7__16_ VDD VSS NOR2_X1 
XU150 A[7] n85 ab_7__17_ VDD VSS NOR2_X1 
XU149 n101 n77 ab_7__1_ VDD VSS NOR2_X1 
XU148 n100 n77 ab_7__2_ VDD VSS NOR2_X1 
XU147 n99 n77 ab_7__3_ VDD VSS NOR2_X1 
XU146 n98 n77 ab_7__4_ VDD VSS NOR2_X1 
XU145 n97 n77 ab_7__5_ VDD VSS NOR2_X1 
XU144 n96 n77 ab_7__6_ VDD VSS NOR2_X1 
XU143 n95 n77 ab_7__7_ VDD VSS NOR2_X1 
XU142 n94 n77 ab_7__8_ VDD VSS NOR2_X1 
XU141 n93 n77 ab_7__9_ VDD VSS NOR2_X1 
XU140 n156 n76 ab_8__0_ VDD VSS NOR2_X1 
XU139 n92 n76 ab_8__10_ VDD VSS NOR2_X1 
XU138 n91 n76 ab_8__11_ VDD VSS NOR2_X1 
XU137 n90 n76 ab_8__12_ VDD VSS NOR2_X1 
XU136 n89 n76 ab_8__13_ VDD VSS NOR2_X1 
XU135 n88 n76 ab_8__14_ VDD VSS NOR2_X1 
XU134 n87 n76 ab_8__15_ VDD VSS NOR2_X1 
XU133 n86 n76 ab_8__16_ VDD VSS NOR2_X1 
XU132 A[8] n85 ab_8__17_ VDD VSS NOR2_X1 
XU131 n101 n76 ab_8__1_ VDD VSS NOR2_X1 
XU130 n100 n76 ab_8__2_ VDD VSS NOR2_X1 
XU129 n99 n76 ab_8__3_ VDD VSS NOR2_X1 
XU128 n98 n76 ab_8__4_ VDD VSS NOR2_X1 
XU127 n97 n76 ab_8__5_ VDD VSS NOR2_X1 
XU126 n96 n76 ab_8__6_ VDD VSS NOR2_X1 
XU125 n95 n76 ab_8__7_ VDD VSS NOR2_X1 
XU124 n94 n76 ab_8__8_ VDD VSS NOR2_X1 
XU123 n93 n76 ab_8__9_ VDD VSS NOR2_X1 
XU122 n75 n156 ab_9__0_ VDD VSS NOR2_X1 
XU121 n75 n92 ab_9__10_ VDD VSS NOR2_X1 
XU120 n75 n91 ab_9__11_ VDD VSS NOR2_X1 
XU305 n95 n71 ab_13__7_ VDD VSS NOR2_X1 
XU304 n94 n71 ab_13__8_ VDD VSS NOR2_X1 
XU303 n93 n71 ab_13__9_ VDD VSS NOR2_X1 
XU302 n156 n35 ab_14__0_ VDD VSS NOR2_X1 
XU301 n92 n35 ab_14__10_ VDD VSS NOR2_X1 
XU300 n91 n35 ab_14__11_ VDD VSS NOR2_X1 
XU299 n90 n35 ab_14__12_ VDD VSS NOR2_X1 
XU298 n89 n35 ab_14__13_ VDD VSS NOR2_X1 
XU297 n88 n35 ab_14__14_ VDD VSS NOR2_X1 
XU296 n87 n35 ab_14__15_ VDD VSS NOR2_X1 
XU295 n86 n35 ab_14__16_ VDD VSS NOR2_X1 
XU294 A[14] n85 ab_14__17_ VDD VSS NOR2_X1 
XU293 n101 n35 ab_14__1_ VDD VSS NOR2_X1 
XU292 n100 n35 ab_14__2_ VDD VSS NOR2_X1 
XU291 n99 n35 ab_14__3_ VDD VSS NOR2_X1 
XU290 n98 n35 ab_14__4_ VDD VSS NOR2_X1 
XU289 n97 n35 ab_14__5_ VDD VSS NOR2_X1 
XU288 n96 n35 ab_14__6_ VDD VSS NOR2_X1 
XU287 n95 n35 ab_14__7_ VDD VSS NOR2_X1 
XU286 n94 n35 ab_14__8_ VDD VSS NOR2_X1 
XU285 n93 n35 ab_14__9_ VDD VSS NOR2_X1 
XU284 B[0] n1 ab_15__0_ VDD VSS NOR2_X1 
XU283 B[10] n1 ab_15__10_ VDD VSS NOR2_X1 
XU282 B[11] n1 ab_15__11_ VDD VSS NOR2_X1 
XU281 B[12] n1 ab_15__12_ VDD VSS NOR2_X1 
XU280 B[13] n1 ab_15__13_ VDD VSS NOR2_X1 
XU279 B[14] n1 ab_15__14_ VDD VSS NOR2_X1 
XU278 B[15] n1 ab_15__15_ VDD VSS NOR2_X1 
XU277 B[16] n1 ab_15__16_ VDD VSS NOR2_X1 
XU276 n85 n1 ab_15__17_ VDD VSS NOR2_X1 
XU275 B[1] n1 ab_15__1_ VDD VSS NOR2_X1 
XU274 B[2] n1 ab_15__2_ VDD VSS NOR2_X1 
XU273 B[3] n1 ab_15__3_ VDD VSS NOR2_X1 
XU272 B[4] n1 ab_15__4_ VDD VSS NOR2_X1 
XU271 B[5] n1 ab_15__5_ VDD VSS NOR2_X1 
XU270 B[6] n1 ab_15__6_ VDD VSS NOR2_X1 
XU269 B[7] n1 ab_15__7_ VDD VSS NOR2_X1 
XU268 B[8] n1 ab_15__8_ VDD VSS NOR2_X1 
XU267 B[9] n1 ab_15__9_ VDD VSS NOR2_X1 
XU266 n156 n83 ab_1__0_ VDD VSS NOR2_X1 
XU265 n92 n83 ab_1__10_ VDD VSS NOR2_X1 
XU264 n91 n83 ab_1__11_ VDD VSS NOR2_X1 
XU263 n90 n83 ab_1__12_ VDD VSS NOR2_X1 
XU262 n89 n83 ab_1__13_ VDD VSS NOR2_X1 
XU261 n88 n83 ab_1__14_ VDD VSS NOR2_X1 
XU260 n87 n83 ab_1__15_ VDD VSS NOR2_X1 
XU259 n86 n83 ab_1__16_ VDD VSS NOR2_X1 
XU258 A[1] n85 ab_1__17_ VDD VSS NOR2_X1 
XU257 n101 n83 ab_1__1_ VDD VSS NOR2_X1 
XU256 n100 n83 ab_1__2_ VDD VSS NOR2_X1 
XU255 n99 n83 ab_1__3_ VDD VSS NOR2_X1 
XU254 n98 n83 ab_1__4_ VDD VSS NOR2_X1 
XU253 n97 n83 ab_1__5_ VDD VSS NOR2_X1 
XU252 n96 n83 ab_1__6_ VDD VSS NOR2_X1 
XU251 n95 n83 ab_1__7_ VDD VSS NOR2_X1 
XU250 n94 n83 ab_1__8_ VDD VSS NOR2_X1 
XU249 n93 n83 ab_1__9_ VDD VSS NOR2_X1 
XU248 n156 n82 ab_2__0_ VDD VSS NOR2_X1 
XU247 n92 n82 ab_2__10_ VDD VSS NOR2_X1 
XU246 n91 n82 ab_2__11_ VDD VSS NOR2_X1 
XU245 n90 n82 ab_2__12_ VDD VSS NOR2_X1 
XU244 n89 n82 ab_2__13_ VDD VSS NOR2_X1 
XU243 n88 n82 ab_2__14_ VDD VSS NOR2_X1 
XU242 n87 n82 ab_2__15_ VDD VSS NOR2_X1 
XU241 n86 n82 ab_2__16_ VDD VSS NOR2_X1 
XU240 A[2] n85 ab_2__17_ VDD VSS NOR2_X1 
XU239 n101 n82 ab_2__1_ VDD VSS NOR2_X1 
XU238 n100 n82 ab_2__2_ VDD VSS NOR2_X1 
XU237 n99 n82 ab_2__3_ VDD VSS NOR2_X1 
XU236 n98 n82 ab_2__4_ VDD VSS NOR2_X1 
XU235 n97 n82 ab_2__5_ VDD VSS NOR2_X1 
XU234 n96 n82 ab_2__6_ VDD VSS NOR2_X1 
XU233 n95 n82 ab_2__7_ VDD VSS NOR2_X1 
XU232 n94 n82 ab_2__8_ VDD VSS NOR2_X1 
XU231 n93 n82 ab_2__9_ VDD VSS NOR2_X1 
XU230 n156 n81 ab_3__0_ VDD VSS NOR2_X1 
XU229 n92 n81 ab_3__10_ VDD VSS NOR2_X1 
XU228 n91 n81 ab_3__11_ VDD VSS NOR2_X1 
XU227 n90 n81 ab_3__12_ VDD VSS NOR2_X1 
XU226 n89 n81 ab_3__13_ VDD VSS NOR2_X1 
XU225 n88 n81 ab_3__14_ VDD VSS NOR2_X1 
XU224 n87 n81 ab_3__15_ VDD VSS NOR2_X1 
XU223 n86 n81 ab_3__16_ VDD VSS NOR2_X1 
XU222 A[3] n85 ab_3__17_ VDD VSS NOR2_X1 
XU221 n101 n81 ab_3__1_ VDD VSS NOR2_X1 
XU220 n100 n81 ab_3__2_ VDD VSS NOR2_X1 
XU219 n99 n81 ab_3__3_ VDD VSS NOR2_X1 
XU218 n98 n81 ab_3__4_ VDD VSS NOR2_X1 
XU217 n97 n81 ab_3__5_ VDD VSS NOR2_X1 
XU216 n96 n81 ab_3__6_ VDD VSS NOR2_X1 
XU215 n95 n81 ab_3__7_ VDD VSS NOR2_X1 
XU214 n94 n81 ab_3__8_ VDD VSS NOR2_X1 
XU213 n93 n81 ab_3__9_ VDD VSS NOR2_X1 
XU392 n156 n84 n157 VDD VSS NOR2_X1 
XU391 n92 n84 ab_0__10_ VDD VSS NOR2_X1 
XU390 n91 n84 ab_0__11_ VDD VSS NOR2_X1 
XU389 n90 n84 ab_0__12_ VDD VSS NOR2_X1 
XU388 n89 n84 ab_0__13_ VDD VSS NOR2_X1 
XU387 n88 n84 ab_0__14_ VDD VSS NOR2_X1 
XU386 n87 n84 ab_0__15_ VDD VSS NOR2_X1 
XU385 n86 n84 ab_0__16_ VDD VSS NOR2_X1 
XU384 A[0] n85 ab_0__17_ VDD VSS NOR2_X1 
XU383 n101 n84 ab_0__1_ VDD VSS NOR2_X1 
XU382 n100 n84 ab_0__2_ VDD VSS NOR2_X1 
XU381 n99 n84 ab_0__3_ VDD VSS NOR2_X1 
XU380 n98 n84 ab_0__4_ VDD VSS NOR2_X1 
XU379 n97 n84 ab_0__5_ VDD VSS NOR2_X1 
XU378 n96 n84 ab_0__6_ VDD VSS NOR2_X1 
XU377 n95 n84 ab_0__7_ VDD VSS NOR2_X1 
XU376 n94 n84 ab_0__8_ VDD VSS NOR2_X1 
XU375 n93 n84 ab_0__9_ VDD VSS NOR2_X1 
XU374 n156 n74 ab_10__0_ VDD VSS NOR2_X1 
XU373 n92 n74 ab_10__10_ VDD VSS NOR2_X1 
XU372 n91 n74 ab_10__11_ VDD VSS NOR2_X1 
XU371 n90 n74 ab_10__12_ VDD VSS NOR2_X1 
XU370 n89 n74 ab_10__13_ VDD VSS NOR2_X1 
XU369 n88 n74 ab_10__14_ VDD VSS NOR2_X1 
XU368 n87 n74 ab_10__15_ VDD VSS NOR2_X1 
XU367 n86 n74 ab_10__16_ VDD VSS NOR2_X1 
XU366 A[10] n85 ab_10__17_ VDD VSS NOR2_X1 
XU365 n101 n74 ab_10__1_ VDD VSS NOR2_X1 
XU364 n100 n74 ab_10__2_ VDD VSS NOR2_X1 
XU363 n99 n74 ab_10__3_ VDD VSS NOR2_X1 
XU362 n98 n74 ab_10__4_ VDD VSS NOR2_X1 
XU361 n97 n74 ab_10__5_ VDD VSS NOR2_X1 
XU360 n96 n74 ab_10__6_ VDD VSS NOR2_X1 
XU359 n95 n74 ab_10__7_ VDD VSS NOR2_X1 
XU358 n94 n74 ab_10__8_ VDD VSS NOR2_X1 
XU357 n93 n74 ab_10__9_ VDD VSS NOR2_X1 
XU356 n156 n73 ab_11__0_ VDD VSS NOR2_X1 
XU355 n92 n73 ab_11__10_ VDD VSS NOR2_X1 
XU354 n91 n73 ab_11__11_ VDD VSS NOR2_X1 
XU353 n90 n73 ab_11__12_ VDD VSS NOR2_X1 
XU352 n89 n73 ab_11__13_ VDD VSS NOR2_X1 
XU351 n88 n73 ab_11__14_ VDD VSS NOR2_X1 
XU350 n87 n73 ab_11__15_ VDD VSS NOR2_X1 
XU349 n86 n73 ab_11__16_ VDD VSS NOR2_X1 
XU348 A[11] n85 ab_11__17_ VDD VSS NOR2_X1 
XU347 n101 n73 ab_11__1_ VDD VSS NOR2_X1 
XU346 n100 n73 ab_11__2_ VDD VSS NOR2_X1 
XU345 n99 n73 ab_11__3_ VDD VSS NOR2_X1 
XU344 n98 n73 ab_11__4_ VDD VSS NOR2_X1 
XU343 n97 n73 ab_11__5_ VDD VSS NOR2_X1 
XU342 n96 n73 ab_11__6_ VDD VSS NOR2_X1 
XU341 n95 n73 ab_11__7_ VDD VSS NOR2_X1 
XU340 n94 n73 ab_11__8_ VDD VSS NOR2_X1 
XU339 n93 n73 ab_11__9_ VDD VSS NOR2_X1 
XU338 n156 n72 ab_12__0_ VDD VSS NOR2_X1 
XU337 n92 n72 ab_12__10_ VDD VSS NOR2_X1 
XU336 n91 n72 ab_12__11_ VDD VSS NOR2_X1 
XU335 n90 n72 ab_12__12_ VDD VSS NOR2_X1 
XU334 n89 n72 ab_12__13_ VDD VSS NOR2_X1 
XU333 n88 n72 ab_12__14_ VDD VSS NOR2_X1 
XU332 n87 n72 ab_12__15_ VDD VSS NOR2_X1 
XU331 n86 n72 ab_12__16_ VDD VSS NOR2_X1 
XU330 A[12] n85 ab_12__17_ VDD VSS NOR2_X1 
XU329 n101 n72 ab_12__1_ VDD VSS NOR2_X1 
XU328 n100 n72 ab_12__2_ VDD VSS NOR2_X1 
XU327 n99 n72 ab_12__3_ VDD VSS NOR2_X1 
XU326 n98 n72 ab_12__4_ VDD VSS NOR2_X1 
XU325 n97 n72 ab_12__5_ VDD VSS NOR2_X1 
XU324 n96 n72 ab_12__6_ VDD VSS NOR2_X1 
XU323 n95 n72 ab_12__7_ VDD VSS NOR2_X1 
XU322 n94 n72 ab_12__8_ VDD VSS NOR2_X1 
XU321 n93 n72 ab_12__9_ VDD VSS NOR2_X1 
XU320 n156 n71 ab_13__0_ VDD VSS NOR2_X1 
XU319 n92 n71 ab_13__10_ VDD VSS NOR2_X1 
XU318 n91 n71 ab_13__11_ VDD VSS NOR2_X1 
XU317 n90 n71 ab_13__12_ VDD VSS NOR2_X1 
XU316 n89 n71 ab_13__13_ VDD VSS NOR2_X1 
XU315 n88 n71 ab_13__14_ VDD VSS NOR2_X1 
XU314 n87 n71 ab_13__15_ VDD VSS NOR2_X1 
XU313 n86 n71 ab_13__16_ VDD VSS NOR2_X1 
XU312 A[13] n85 ab_13__17_ VDD VSS NOR2_X1 
XU311 n101 n71 ab_13__1_ VDD VSS NOR2_X1 
XU310 n100 n71 ab_13__2_ VDD VSS NOR2_X1 
XU309 n99 n71 ab_13__3_ VDD VSS NOR2_X1 
XU308 n98 n71 ab_13__4_ VDD VSS NOR2_X1 
XU307 n97 n71 ab_13__5_ VDD VSS NOR2_X1 
XU306 n96 n71 ab_13__6_ VDD VSS NOR2_X1 
XU104 n119 PRODUCT[14] VDD VSS BUF_X1 
XU393 n127 PRODUCT[10] VDD VSS BUF_X1 
XU394 n129 PRODUCT[9] VDD VSS BUF_X1 
XU395 n134 PRODUCT[7] VDD VSS BUF_X1 
XU396 n136 PRODUCT[6] VDD VSS BUF_X1 
XU397 n138 PRODUCT[5] VDD VSS BUF_X1 
XU398 n139 PRODUCT[4] VDD VSS BUF_X1 
XU399 n143 PRODUCT[3] VDD VSS BUF_X1 
XU400 n144 PRODUCT[2] VDD VSS BUF_X1 
XU401 n148 PRODUCT[1] VDD VSS BUF_X1 
XU402 n152 PRODUCT[0] VDD VSS BUF_X1 
XU403 n102 n155 VDD VSS INV_X1 
XU404 n145 n146 VDD VSS INV_X1 
XU405 n137 n138 VDD VSS INV_X16 
XU406 n140 n141 VDD VSS INV_X1 
XU407 n131 n132 VDD VSS INV_X1 
XU408 n118 n119 VDD VSS INV_X16 
XU409 n117 n114 VDD VSS INV_X1 
XU410 n114 PRODUCT[15] VDD VSS INV_X32 
XU411 n69 n116 VDD VSS INV_X1 
XU412 n116 n117 VDD VSS INV_X32 
XU413 A1_12_ n118 VDD VSS INV_X32 
XU414 A1_11_ n120 VDD VSS INV_X32 
XU415 n120 PRODUCT[13] VDD VSS INV_X32 
XU416 A1_10_ n122 VDD VSS INV_X32 
XU417 n122 PRODUCT[12] VDD VSS INV_X32 
XU418 A1_9_ n124 VDD VSS INV_X32 
XU419 n124 n125 VDD VSS INV_X32 
XU420 A1_8_ n126 VDD VSS INV_X32 
XU421 n126 n127 VDD VSS INV_X16 
XU422 A1_7_ n128 VDD VSS INV_X32 
XU423 n128 n129 VDD VSS INV_X32 
XU424 n132 n130 VDD VSS BUF_X1 
XU425 A1_6_ n131 VDD VSS INV_X32 
XU426 A1_5_ n133 VDD VSS INV_X32 
XU427 n133 n134 VDD VSS INV_X32 
XU428 A1_4_ n135 VDD VSS INV_X32 
XU429 n135 n136 VDD VSS INV_X32 
XU430 A1_3_ n137 VDD VSS INV_X32 
XU431 n141 n139 VDD VSS BUF_X1 
XU432 A1_2_ n140 VDD VSS INV_X32 
XU433 A1_1_ n142 VDD VSS INV_X32 
XU434 n142 n143 VDD VSS INV_X32 
XU435 n146 n144 VDD VSS BUF_X1 
XU436 A1_0_ n145 VDD VSS INV_X32 
XU437 n150 n147 VDD VSS INV_X1 
XU438 n147 n148 VDD VSS INV_X16 
XU439 n158 n149 VDD VSS INV_X1 
XU440 n149 n150 VDD VSS INV_X32 
XU441 n154 n151 VDD VSS INV_X1 
XU442 n151 n152 VDD VSS INV_X32 
XU443 n157 n153 VDD VSS INV_X1 
XU444 n153 n154 VDD VSS INV_X32 
XU445 n155 n156 VDD VSS INV_X1 
XU461 n125 PRODUCT[11] VDD VSS BUF_X1 
XU462 n130 PRODUCT[8] VDD VSS BUF_X1 
XFS_1 VSS SYNOPSYS_UNCONNECTED_94 VDD VSS PRODUCT[33] PRODUCT[32] PRODUCT[31] PRODUCT[30] 
+ PRODUCT[29] PRODUCT[28] PRODUCT[27] PRODUCT[26] PRODUCT[25] PRODUCT[24] PRODUCT[23] 
+ PRODUCT[22] PRODUCT[21] PRODUCT[20] PRODUCT[19] PRODUCT[18] PRODUCT[17] PRODUCT[16] 
+ n49 n61 n60 n59 n58 n57 n56 n55 n54 n53 n52 n51 n50 n41 n40 A2_16_ n39 n68 VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS n70 n48 n67 n47 n66 n46 n65 
+ n45 n64 n44 n63 n43 n62 n37 n42 n36 A1_15_ n38 PRODUCT[15] PRODUCT[14] PRODUCT[13] 
+ PRODUCT[12] PRODUCT[11] PRODUCT[10] PRODUCT[9] PRODUCT[8] PRODUCT[7] PRODUCT[6] 
+ PRODUCT[5] PRODUCT[4] PRODUCT[3] PRODUCT[2] gng_smul_16_18_sadd_37_DW01_add_1 
.ENDS

.SUBCKT gng_smul_16_18_sadd_37 p[37] p[36] p[35] p[34] p[33] p[32] p[31] p[30] p[29] 
+ p[28] p[27] p[26] p[25] p[24] p[23] p[22] p[21] p[20] p[19] p[18] p[17] p[16] 
+ p[15] p[14] p[13] p[12] p[11] p[10] p[9] p[8] p[7] p[6] p[5] p[4] p[3] p[2] p[1] 
+ p[0] clk VDD VSS c[36] c[35] c[34] c[33] c[32] c[31] c[30] c[29] c[28] c[27] c[26] 
+ c[25] c[24] c[23] c[22] c[21] c[20] c[19] c[18] c[17] c[16] c[15] c[14] c[13] 
+ c[12] c[11] c[10] c[9] c[8] c[7] c[6] c[5] c[4] c[3] c[2] c[1] c[0] b[17] b[16] 
+ b[15] b[14] b[13] b[12] b[11] b[10] b[9] b[8] b[7] b[6] b[5] b[4] b[3] b[2] b[1] 
+ b[0] a[15] a[14] a[13] a[12] a[11] a[10] a[9] a[8] a[7] a[6] a[5] a[4] a[3] a[2] 
+ a[1] a[0] 
XLOGIC0_X1_U1 LOGIC0_X1_U1_net VDD VSS LOGIC0_X1 
XLOGIC0_X1_U2 LOGIC0_X1_U2_net VDD VSS LOGIC0_X1 
XLOGIC0_X1_U3 LOGIC0_X1_U3_net VDD VSS LOGIC0_X1 
XLOGIC0_X1_U4 LOGIC0_X1_U4_net VDD VSS LOGIC0_X1 
Xprod_reg_30_ N301 n2_G3B1I6 prod[30] SYNOPSYS_UNCONNECTED_219 VDD VSS DFF_X1 
Xprod_reg_31_ N310 n2_G3B1I6 prod[31] SYNOPSYS_UNCONNECTED_218 VDD VSS DFF_X1 
Xprod_reg_32_ N320 n2_G3B1I2 prod[32] SYNOPSYS_UNCONNECTED_217 VDD VSS DFF_X1 
Xprod_reg_33_ N33 n2_G3B1I2 prod[33] SYNOPSYS_UNCONNECTED_216 VDD VSS DFF_X1 
Xc_reg_reg_0_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[0] SYNOPSYS_UNCONNECTED_215 VDD VSS DFF_X1 
Xc_reg_reg_1_ LOGIC0_X1_U4_net n3 c_reg[1] SYNOPSYS_UNCONNECTED_214 VDD VSS DFF_X1 
Xc_reg_reg_2_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[2] SYNOPSYS_UNCONNECTED_213 VDD VSS DFF_X1 
Xc_reg_reg_3_ LOGIC0_X1_U4_net n3 c_reg[3] SYNOPSYS_UNCONNECTED_212 VDD VSS DFF_X1 
Xc_reg_reg_4_ LOGIC0_X1_U4_net n3 c_reg[4] SYNOPSYS_UNCONNECTED_211 VDD VSS DFF_X1 
Xc_reg_reg_5_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[5] SYNOPSYS_UNCONNECTED_210 VDD VSS DFF_X1 
Xc_reg_reg_6_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[6] SYNOPSYS_UNCONNECTED_209 VDD VSS DFF_X1 
Xc_reg_reg_7_ LOGIC0_X1_U4_net n3_G3B1I4 c_reg[7] SYNOPSYS_UNCONNECTED_208 VDD VSS DFF_X1 
Xc_reg_reg_8_ LOGIC0_X1_U3_net n3_G3B1I4 c_reg[8] SYNOPSYS_UNCONNECTED_207 VDD VSS DFF_X1 
Xc_reg_reg_9_ LOGIC0_X1_U4_net n3_G3B1I4 c_reg[9] SYNOPSYS_UNCONNECTED_206 VDD VSS DFF_X1 
Xc_reg_reg_10_ LOGIC0_X1_U4_net n3_G3B1I3 c_reg[10] SYNOPSYS_UNCONNECTED_205 VDD 
+ VSS DFF_X1 
Xc_reg_reg_11_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[11] SYNOPSYS_UNCONNECTED_204 VDD 
+ VSS DFF_X1 
Xc_reg_reg_12_ LOGIC0_X1_U1_net n3_G3B1I5 c_reg[12] SYNOPSYS_UNCONNECTED_203 VDD 
+ VSS DFF_X1 
Xc_reg_reg_13_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[13] SYNOPSYS_UNCONNECTED_202 VDD 
+ VSS DFF_X1 
Xc_reg_reg_14_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[14] SYNOPSYS_UNCONNECTED_201 VDD 
+ VSS DFF_X1 
Xc_reg_reg_15_ LOGIC0_X1_U1_net n3_G3B1I2 c_reg[15] SYNOPSYS_UNCONNECTED_200 VDD 
+ VSS DFF_X1 
Xc_reg_reg_16_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[16] SYNOPSYS_UNCONNECTED_199 VDD 
+ VSS DFF_X1 
Xc_reg_reg_17_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[17] SYNOPSYS_UNCONNECTED_198 VDD 
+ VSS DFF_X1 
Xc_reg_reg_18_ LOGIC0_X1_U2_net n1_G3B1I5 c_reg[18] SYNOPSYS_UNCONNECTED_197 VDD 
+ VSS DFF_X1 
Xc_reg_reg_19_ c[19] n1_G3B1I6 c_reg[19] SYNOPSYS_UNCONNECTED_196 VDD VSS DFF_X1 
Xc_reg_reg_20_ c[20] n1_G3B1I3 c_reg[20] SYNOPSYS_UNCONNECTED_195 VDD VSS DFF_X1 
Xc_reg_reg_21_ c[21] n1_G3B1I3 c_reg[21] SYNOPSYS_UNCONNECTED_194 VDD VSS DFF_X1 
Xc_reg_reg_22_ c[22] n1_G3B1I3 c_reg[22] SYNOPSYS_UNCONNECTED_193 VDD VSS DFF_X1 
Xc_reg_reg_23_ c[23] n1_G3B1I3 c_reg[23] SYNOPSYS_UNCONNECTED_192 VDD VSS DFF_X1 
Xc_reg_reg_24_ c[24] n2_G3B1I3 c_reg[24] SYNOPSYS_UNCONNECTED_191 VDD VSS DFF_X1 
Xc_reg_reg_25_ c[25] n2_G3B1I3 c_reg[25] SYNOPSYS_UNCONNECTED_190 VDD VSS DFF_X1 
Xc_reg_reg_26_ c[26] n2_G3B1I3 c_reg[26] SYNOPSYS_UNCONNECTED_189 VDD VSS DFF_X1 
Xc_reg_reg_27_ c[27] n2_G3B1I3 c_reg[27] SYNOPSYS_UNCONNECTED_188 VDD VSS DFF_X1 
Xc_reg_reg_28_ c[28] n2_G3B1I3 c_reg[28] SYNOPSYS_UNCONNECTED_187 VDD VSS DFF_X1 
Xc_reg_reg_29_ c[29] n2_G3B1I3 c_reg[29] SYNOPSYS_UNCONNECTED_186 VDD VSS DFF_X1 
Xc_reg_reg_30_ c[30] n2_G3B1I3 c_reg[30] SYNOPSYS_UNCONNECTED_185 VDD VSS DFF_X1 
Xc_reg_reg_31_ c[31] n2_G3B1I4 c_reg[31] SYNOPSYS_UNCONNECTED_184 VDD VSS DFF_X1 
Xc_reg_reg_32_ c[32] n2_G3B1I4 c_reg[32] SYNOPSYS_UNCONNECTED_183 VDD VSS DFF_X1 
Xc_reg_reg_33_ c[33] n2_G3B1I4 c_reg[33] SYNOPSYS_UNCONNECTED_182 VDD VSS DFF_X1 
Xc_reg_reg_34_ c[34] n2_G3B1I2 c_reg[34] SYNOPSYS_UNCONNECTED_181 VDD VSS DFF_X1 
Xc_reg_reg_35_ c[35] n2_G3B1I2 c_reg[35] SYNOPSYS_UNCONNECTED_180 VDD VSS DFF_X1 
Xc_reg_reg_36_ c[36] n2_G3B1I2 c_reg[36] SYNOPSYS_UNCONNECTED_179 VDD VSS DFF_X1 
Xb_reg_reg_0_ b[0] n2_G3B1I1 b_reg[0] SYNOPSYS_UNCONNECTED_178 VDD VSS DFF_X1 
Xb_reg_reg_1_ b[1] n2_G3B1I1 b_reg[1] SYNOPSYS_UNCONNECTED_177 VDD VSS DFF_X1 
Xb_reg_reg_2_ b[2] n1_G3B1I6 b_reg[2] SYNOPSYS_UNCONNECTED_176 VDD VSS DFF_X1 
Xb_reg_reg_3_ b[3] n1_G3B1I6 b_reg[3] SYNOPSYS_UNCONNECTED_175 VDD VSS DFF_X1 
Xb_reg_reg_4_ b[4] n1_G3B1I2 b_reg[4] SYNOPSYS_UNCONNECTED_174 VDD VSS DFF_X1 
Xb_reg_reg_5_ b[5] n1_G3B1I2 b_reg[5] SYNOPSYS_UNCONNECTED_173 VDD VSS DFF_X1 
Xb_reg_reg_6_ b[6] n1_G3B1I2 b_reg[6] SYNOPSYS_UNCONNECTED_172 VDD VSS DFF_X1 
Xb_reg_reg_7_ b[7] n1_G3B1I3 b_reg[7] SYNOPSYS_UNCONNECTED_171 VDD VSS DFF_X1 
Xb_reg_reg_8_ b[8] n1_G3B1I4 b_reg[8] SYNOPSYS_UNCONNECTED_170 VDD VSS DFF_X1 
Xb_reg_reg_9_ b[9] n1_G3B1I4 b_reg[9] SYNOPSYS_UNCONNECTED_169 VDD VSS DFF_X1 
Xb_reg_reg_10_ b[10] n2_G3B1I1 b_reg[10] SYNOPSYS_UNCONNECTED_168 VDD VSS DFF_X1 
Xb_reg_reg_11_ b[11] n2_G3B1I6 b_reg[11] SYNOPSYS_UNCONNECTED_167 VDD VSS DFF_X1 
Xb_reg_reg_12_ b[12] n2_G3B1I1 b_reg[12] SYNOPSYS_UNCONNECTED_166 VDD VSS DFF_X1 
Xb_reg_reg_13_ b[13] n2_G3B1I6 b_reg[13] SYNOPSYS_UNCONNECTED_165 VDD VSS DFF_X1 
Xb_reg_reg_14_ b[14] n2_G3B1I1 b_reg[14] SYNOPSYS_UNCONNECTED_164 VDD VSS DFF_X1 
Xb_reg_reg_15_ b[15] n2_G3B1I1 b_reg[15] SYNOPSYS_UNCONNECTED_163 VDD VSS DFF_X1 
Xb_reg_reg_16_ b[16] n2_G3B1I1 b_reg[16] SYNOPSYS_UNCONNECTED_162 VDD VSS DFF_X1 
Xb_reg_reg_17_ LOGIC0_X1_U2_net n1_G3B1I2 b_reg[17] SYNOPSYS_UNCONNECTED_161 VDD 
+ VSS DFF_X1 
Xa_reg_reg_0_ a[0] n1_G3B1I6 a_reg[0] SYNOPSYS_UNCONNECTED_160 VDD VSS DFF_X1 
Xa_reg_reg_1_ a[1] n1_G3B1I6 a_reg[1] SYNOPSYS_UNCONNECTED_159 VDD VSS DFF_X1 
Xa_reg_reg_2_ a[2] n1_G3B1I2 a_reg[2] SYNOPSYS_UNCONNECTED_158 VDD VSS DFF_X1 
Xa_reg_reg_3_ a[3] n1_G3B1I6 a_reg[3] SYNOPSYS_UNCONNECTED_157 VDD VSS DFF_X1 
Xa_reg_reg_4_ a[4] n1_G3B1I1 a_reg[4] SYNOPSYS_UNCONNECTED_156 VDD VSS DFF_X1 
Xa_reg_reg_5_ a[5] n1_G3B1I2 a_reg[5] SYNOPSYS_UNCONNECTED_155 VDD VSS DFF_X1 
Xa_reg_reg_6_ a[6] n1_G3B1I1 a_reg[6] SYNOPSYS_UNCONNECTED_154 VDD VSS DFF_X1 
Xa_reg_reg_7_ a[7] n1_G3B1I1 a_reg[7] SYNOPSYS_UNCONNECTED_153 VDD VSS DFF_X1 
Xa_reg_reg_8_ a[8] n1_G3B1I1 a_reg[8] SYNOPSYS_UNCONNECTED_152 VDD VSS DFF_X1 
Xa_reg_reg_9_ a[9] n2 a_reg[9] SYNOPSYS_UNCONNECTED_151 VDD VSS DFF_X1 
Xa_reg_reg_10_ a[10] n1_G3B1I4 a_reg[10] SYNOPSYS_UNCONNECTED_150 VDD VSS DFF_X1 
Xa_reg_reg_11_ a[11] n1_G3B1I4 a_reg[11] SYNOPSYS_UNCONNECTED_149 VDD VSS DFF_X1 
Xa_reg_reg_12_ a[12] n1_G3B1I4 a_reg[12] SYNOPSYS_UNCONNECTED_148 VDD VSS DFF_X1 
Xa_reg_reg_13_ a[13] n1_G3B1I4 a_reg[13] SYNOPSYS_UNCONNECTED_147 VDD VSS DFF_X1 
Xa_reg_reg_14_ a[14] n1_G3B1I4 a_reg[14] SYNOPSYS_UNCONNECTED_146 VDD VSS DFF_X1 
Xa_reg_reg_15_ LOGIC0_X1_U2_net n1_G3B1I1 a_reg[15] SYNOPSYS_UNCONNECTED_145 VDD 
+ VSS DFF_X1 
Xresult_reg_20_ sum[20] n1_G3B1I3 n119 SYNOPSYS_UNCONNECTED_144 VDD VSS DFF_X1 
Xresult_reg_21_ sum[21] n1_G3B1I3 n120 SYNOPSYS_UNCONNECTED_143 VDD VSS DFF_X1 
Xresult_reg_22_ sum[22] n1_G3B1I4 n121 SYNOPSYS_UNCONNECTED_142 VDD VSS DFF_X1 
Xresult_reg_23_ sum[23] n1_G3B1I4 n122 SYNOPSYS_UNCONNECTED_141 VDD VSS DFF_X1 
Xresult_reg_24_ sum[24] n2_G3B1I2 n123 SYNOPSYS_UNCONNECTED_140 VDD VSS DFF_X1 
Xresult_reg_25_ n124 n2_G3B1I3 n111 SYNOPSYS_UNCONNECTED_139 VDD VSS DFF_X1 
Xresult_reg_26_ sum[26] n2_G3B1I5 n112 SYNOPSYS_UNCONNECTED_138 VDD VSS DFF_X1 
Xresult_reg_27_ sum[27] n2_G3B1I5 n113 SYNOPSYS_UNCONNECTED_137 VDD VSS DFF_X1 
Xresult_reg_28_ sum[28] n2_G3B1I5 n114 SYNOPSYS_UNCONNECTED_136 VDD VSS DFF_X1 
Xresult_reg_29_ sum[29] n2_G3B1I5 n115 SYNOPSYS_UNCONNECTED_135 VDD VSS DFF_X1 
Xresult_reg_30_ sum[30] n2_G3B1I5 n116 SYNOPSYS_UNCONNECTED_134 VDD VSS DFF_X1 
Xresult_reg_31_ sum[31] n2_G3B1I4 n117 SYNOPSYS_UNCONNECTED_133 VDD VSS DFF_X1 
Xresult_reg_32_ sum[32] n2_G3B1I4 n118 SYNOPSYS_UNCONNECTED_132 VDD VSS DFF_X1 
Xresult_reg_33_ sum[33] n2_G3B1I4 n106 SYNOPSYS_UNCONNECTED_131 VDD VSS DFF_X1 
Xresult_reg_34_ sum[34] n2_G3B1I4 n107 SYNOPSYS_UNCONNECTED_130 VDD VSS DFF_X1 
Xresult_reg_35_ sum[35] n2_G3B1I2 n108 SYNOPSYS_UNCONNECTED_129 VDD VSS DFF_X1 
Xresult_reg_36_ sum[36] n2_G3B1I2 n109 SYNOPSYS_UNCONNECTED_128 VDD VSS DFF_X1 
Xresult_reg_37_ sum[37] n2_G3B1I6 n110 SYNOPSYS_UNCONNECTED_127 VDD VSS DFF_X1 
Xprod_reg_0_ N0 n3_G3B1I5 prod[0] SYNOPSYS_UNCONNECTED_126 VDD VSS DFF_X1 
Xprod_reg_1_ N1000 n3_G3B1I5 prod[1] SYNOPSYS_UNCONNECTED_125 VDD VSS DFF_X1 
Xprod_reg_2_ N200 n3_G3B1I5 prod[2] SYNOPSYS_UNCONNECTED_124 VDD VSS DFF_X1 
Xprod_reg_3_ N300 n3_G3B1I5 prod[3] SYNOPSYS_UNCONNECTED_123 VDD VSS DFF_X1 
Xprod_reg_4_ N4 n3_G3B1I5 prod[4] SYNOPSYS_UNCONNECTED_122 VDD VSS DFF_X1 
Xprod_reg_5_ N5 n3_G3B1I3 prod[5] SYNOPSYS_UNCONNECTED_121 VDD VSS DFF_X1 
Xprod_reg_6_ N6 n3_G3B1I3 prod[6] SYNOPSYS_UNCONNECTED_120 VDD VSS DFF_X1 
Xprod_reg_7_ N7 n3_G3B1I4 prod[7] SYNOPSYS_UNCONNECTED_119 VDD VSS DFF_X1 
Xprod_reg_8_ N8 n3_G3B1I4 prod[8] SYNOPSYS_UNCONNECTED_118 VDD VSS DFF_X1 
Xprod_reg_9_ N9 n3_G3B1I4 prod[9] SYNOPSYS_UNCONNECTED_117 VDD VSS DFF_X1 
Xprod_reg_10_ N102 n3_G3B1I3 prod[10] SYNOPSYS_UNCONNECTED_116 VDD VSS DFF_X1 
Xprod_reg_11_ N11 n3_G3B1I2 prod[11] SYNOPSYS_UNCONNECTED_115 VDD VSS DFF_X1 
Xprod_reg_12_ N12 n3_G3B1I2 prod[12] SYNOPSYS_UNCONNECTED_114 VDD VSS DFF_X1 
Xprod_reg_13_ N13 n3_G3B1I2 prod[13] SYNOPSYS_UNCONNECTED_113 VDD VSS DFF_X1 
Xprod_reg_14_ N14 n3_G3B1I2 prod[14] SYNOPSYS_UNCONNECTED_112 VDD VSS DFF_X1 
Xprod_reg_15_ N15 n3_G3B1I2 prod[15] SYNOPSYS_UNCONNECTED_111 VDD VSS DFF_X1 
Xprod_reg_16_ N16 n1_G3B1I5 prod[16] SYNOPSYS_UNCONNECTED_110 VDD VSS DFF_X1 
Xprod_reg_17_ N17 n1_G3B1I5 prod[17] SYNOPSYS_UNCONNECTED_109 VDD VSS DFF_X1 
Xprod_reg_18_ N18 n1_G3B1I5 prod[18] SYNOPSYS_UNCONNECTED_108 VDD VSS DFF_X1 
Xprod_reg_19_ N19 n1_G3B1I6 prod[19] SYNOPSYS_UNCONNECTED_107 VDD VSS DFF_X1 
Xprod_reg_20_ N201 n1_G3B1I6 prod[20] SYNOPSYS_UNCONNECTED_106 VDD VSS DFF_X1 
Xprod_reg_21_ N21 n1_G3B1I3 prod[21] SYNOPSYS_UNCONNECTED_105 VDD VSS DFF_X1 
Xprod_reg_22_ N22 n1_G3B1I3 prod[22] SYNOPSYS_UNCONNECTED_104 VDD VSS DFF_X1 
Xprod_reg_23_ N23 n1_G3B1I4 prod[23] SYNOPSYS_UNCONNECTED_103 VDD VSS DFF_X1 
Xprod_reg_24_ N24 n2_G3B1I1 prod[24] SYNOPSYS_UNCONNECTED_102 VDD VSS DFF_X1 
Xprod_reg_25_ N25 n2_G3B1I6 prod[25] SYNOPSYS_UNCONNECTED_101 VDD VSS DFF_X1 
Xprod_reg_26_ N26 n2_G3B1I6 prod[26] SYNOPSYS_UNCONNECTED_100 VDD VSS DFF_X1 
Xprod_reg_27_ N27 n2_G3B1I6 prod[27] SYNOPSYS_UNCONNECTED_99 VDD VSS DFF_X1 
Xprod_reg_28_ N28 n2_G3B1I6 prod[28] SYNOPSYS_UNCONNECTED_98 VDD VSS DFF_X1 
Xprod_reg_29_ N290 n2_G3B1I6 prod[29] SYNOPSYS_UNCONNECTED_97 VDD VSS DFF_X1 
XU1 clk n1 VDD VSS BUF_X32 
XU2 clk n2 VDD VSS BUF_X32 
XU3 clk n3 VDD VSS BUF_X32 
XCLKBUF_X1_G3B1I61 n1 n1_G3B1I6 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I52 n1 n1_G3B1I5 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I32 n1 n1_G3B1I3 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I22 n1 n1_G3B1I2 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I12 n1 n1_G3B1I1 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I5 n3 n3_G3B1I5 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I4 n3 n3_G3B1I4 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I3 n3 n3_G3B1I3 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I2 n3 n3_G3B1I2 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I6 n2 n2_G3B1I6 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I51 n2 n2_G3B1I5 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I41 n2 n2_G3B1I4 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I31 n2 n2_G3B1I3 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I21 n2 n2_G3B1I2 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I11 n2 n2_G3B1I1 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I42 n1 n1_G3B1I4 VDD VSS CLKBUF_X2 
XU4 n31 n330 VDD VSS INV_X16 
XU5 b_reg[17] n29 VDD VSS INV_X16 
XU6 a_reg[15] n32 VDD VSS INV_X1 
XU7 n29 n302 VDD VSS INV_X1 
XU8 n32 n31 VDD VSS CLKBUF_X1 
XU9 n110 n34 VDD VSS CLKBUF_X1 
XU10 n36 n35 VDD VSS CLKBUF_X1 
XU11 n34 n36 VDD VSS INV_X32 
XU12 n35 p[37] VDD VSS INV_X32 
XU13 n109 n38 VDD VSS CLKBUF_X1 
XU14 n40 n39 VDD VSS CLKBUF_X1 
XU15 n38 n40 VDD VSS INV_X32 
XU16 n39 p[36] VDD VSS INV_X32 
XU17 n108 n42 VDD VSS CLKBUF_X1 
XU18 n44 n43 VDD VSS CLKBUF_X1 
XU19 n42 n44 VDD VSS INV_X32 
XU20 n43 p[35] VDD VSS INV_X32 
XU21 n107 n46 VDD VSS CLKBUF_X1 
XU22 n48 n47 VDD VSS CLKBUF_X1 
XU23 n46 n48 VDD VSS INV_X32 
XU24 n47 p[34] VDD VSS INV_X32 
XU25 n106 n50 VDD VSS CLKBUF_X1 
XU26 n52 n51 VDD VSS CLKBUF_X1 
XU27 n50 n52 VDD VSS INV_X32 
XU28 n51 p[33] VDD VSS INV_X32 
XU29 n118 n54 VDD VSS CLKBUF_X1 
XU30 n56 n55 VDD VSS CLKBUF_X1 
XU31 n54 n56 VDD VSS INV_X32 
XU32 n55 p[32] VDD VSS INV_X32 
XU33 n117 n58 VDD VSS CLKBUF_X1 
XU34 n60 n59 VDD VSS CLKBUF_X1 
XU35 n58 n60 VDD VSS INV_X32 
XU36 n59 p[31] VDD VSS INV_X32 
XU37 n116 n62 VDD VSS CLKBUF_X1 
XU38 n64 n63 VDD VSS CLKBUF_X1 
XU39 n62 n64 VDD VSS INV_X32 
XU40 n63 p[30] VDD VSS INV_X32 
XU41 n115 n66 VDD VSS CLKBUF_X1 
XU42 n68 n67 VDD VSS CLKBUF_X1 
XU43 n66 n68 VDD VSS INV_X32 
XU44 n67 p[29] VDD VSS INV_X32 
XU45 n114 n70 VDD VSS CLKBUF_X1 
XU46 n72 n71 VDD VSS CLKBUF_X1 
XU47 n70 n72 VDD VSS INV_X32 
XU48 n71 p[28] VDD VSS INV_X32 
XU49 n113 n74 VDD VSS CLKBUF_X1 
XU50 n76 n75 VDD VSS CLKBUF_X1 
XU51 n74 n76 VDD VSS INV_X32 
XU52 n75 p[27] VDD VSS INV_X32 
XU53 n112 n78 VDD VSS CLKBUF_X1 
XU54 n80 n79 VDD VSS CLKBUF_X1 
XU55 n78 n80 VDD VSS INV_X32 
XU56 n79 p[26] VDD VSS INV_X32 
XU57 n111 n82 VDD VSS CLKBUF_X1 
XU58 n84 n83 VDD VSS CLKBUF_X1 
XU59 n82 n84 VDD VSS INV_X32 
XU60 n83 p[25] VDD VSS INV_X32 
XU61 n123 n86 VDD VSS CLKBUF_X1 
XU62 n88 n87 VDD VSS CLKBUF_X1 
XU63 n86 n88 VDD VSS INV_X32 
XU64 n87 p[24] VDD VSS INV_X32 
XU65 n122 n90 VDD VSS CLKBUF_X1 
XU66 n92 n91 VDD VSS CLKBUF_X1 
XU67 n90 n92 VDD VSS INV_X32 
XU68 n91 p[23] VDD VSS INV_X32 
XU69 n121 n94 VDD VSS CLKBUF_X1 
XU70 n96 n95 VDD VSS CLKBUF_X1 
XU71 n94 n96 VDD VSS INV_X32 
XU72 n95 p[22] VDD VSS INV_X32 
XU73 n101 p[21] VDD VSS BUF_X1 
XU74 n100 n99 VDD VSS CLKBUF_X1 
XU75 n120 n100 VDD VSS INV_X32 
XU76 n99 n101 VDD VSS INV_X32 
XU77 n105 p[20] VDD VSS BUF_X1 
XU78 n104 n103 VDD VSS CLKBUF_X1 
XU79 n119 n104 VDD VSS INV_X32 
XU80 n103 n105 VDD VSS INV_X32 
XU81 sum[25] n124 VDD VSS BUF_X1 
Xadd_69 sum[37] sum[36] sum[35] sum[34] sum[33] sum[32] sum[31] sum[30] sum[29] 
+ sum[28] sum[27] sum[26] sum[25] sum[24] sum[23] sum[22] sum[21] sum[20] sum[19] 
+ sum[18] sum[17] sum[16] sum[15] sum[14] sum[13] sum[12] sum[11] sum[10] sum[9] 
+ sum[8] sum[7] sum[6] sum[5] sum[4] sum[3] sum[2] sum[1] sum[0] VSS SYNOPSYS_UNCONNECTED_96 
+ VDD VSS prod[33] prod[33] prod[33] prod[33] prod[33] prod[32] prod[31] prod[30] 
+ prod[29] prod[28] prod[27] prod[26] prod[25] prod[24] prod[23] prod[22] prod[21] 
+ prod[20] prod[19] prod[18] prod[17] prod[16] prod[15] prod[14] prod[13] prod[12] 
+ prod[11] prod[10] prod[9] prod[8] prod[7] prod[6] prod[5] prod[4] prod[3] prod[2] 
+ prod[1] prod[0] c_reg[36] c_reg[36] c_reg[35] c_reg[34] c_reg[33] c_reg[32] c_reg[31] 
+ c_reg[30] c_reg[29] c_reg[28] c_reg[27] c_reg[26] c_reg[25] c_reg[24] c_reg[23] 
+ c_reg[22] c_reg[21] c_reg[20] c_reg[19] c_reg[18] c_reg[17] c_reg[16] c_reg[15] 
+ c_reg[14] c_reg[13] c_reg[12] c_reg[11] c_reg[10] c_reg[9] c_reg[8] c_reg[7] c_reg[6] 
+ c_reg[5] c_reg[4] c_reg[3] c_reg[2] c_reg[1] c_reg[0] gng_smul_16_18_sadd_37_DW01_add_0 
Xmult_66 N33 N320 N310 N301 N290 N28 N27 N26 N25 N24 N23 N22 N21 N201 N19 N18 N17 
+ N16 N15 N14 N13 N12 N11 N102 N9 N8 N7 N6 N5 N4 N300 N200 N1000 N0 VDD VDD VSS 
+ n302 b_reg[16] b_reg[15] b_reg[14] b_reg[13] b_reg[12] b_reg[11] b_reg[10] b_reg[9] 
+ b_reg[8] b_reg[7] b_reg[6] b_reg[5] b_reg[4] b_reg[3] b_reg[2] b_reg[1] b_reg[0] 
+ n330 a_reg[14] a_reg[13] a_reg[12] a_reg[11] a_reg[10] a_reg[9] a_reg[8] a_reg[7] 
+ a_reg[6] a_reg[5] a_reg[4] a_reg[3] a_reg[2] a_reg[1] a_reg[0] gng_smul_16_18_sadd_37_DW02_mult_0 
.ENDS

.SUBCKT gng_smul_16_18 p[33] p[32] p[31] p[30] p[29] p[28] p[27] p[26] p[25] p[24] 
+ p[23] p[22] p[21] p[20] p[19] p[18] p[17] p[16] p[15] p[14] p[13] p[12] p[11] 
+ p[10] p[9] p[8] p[7] p[6] p[5] p[4] p[3] p[2] p[1] p[0] clk VDD VSS b[17] b[16] 
+ b[15] b[14] b[13] b[12] b[11] b[10] b[9] b[8] b[7] b[6] b[5] b[4] b[3] b[2] b[1] 
+ b[0] a[15] a[14] a[13] a[12] a[11] a[10] a[9] a[8] a[7] a[6] a[5] a[4] a[3] a[2] 
+ a[1] a[0] 
XLOGIC0_X1_U0 LOGIC0_X1_U0_net VDD VSS LOGIC0_X1 
Xprod_reg_19_ N19 n1_G3B1I4 p[19] SYNOPSYS_UNCONNECTED_93 VDD VSS DFF_X1 
Xprod_reg_20_ N20 n1_G3B1I4 p[20] SYNOPSYS_UNCONNECTED_92 VDD VSS DFF_X1 
Xprod_reg_21_ N21 n1_G3B1I3 p[21] SYNOPSYS_UNCONNECTED_91 VDD VSS DFF_X1 
Xprod_reg_22_ N22 n1_G3B1I2 p[22] SYNOPSYS_UNCONNECTED_90 VDD VSS DFF_X1 
Xprod_reg_23_ N23 n1_G3B1I2 p[23] SYNOPSYS_UNCONNECTED_89 VDD VSS DFF_X1 
Xprod_reg_24_ N24 n1_G3B1I2 p[24] SYNOPSYS_UNCONNECTED_88 VDD VSS DFF_X1 
Xprod_reg_25_ N25 n1_G3B1I2 p[25] SYNOPSYS_UNCONNECTED_87 VDD VSS DFF_X1 
Xprod_reg_26_ N26 n1_G3B1I3 p[26] SYNOPSYS_UNCONNECTED_86 VDD VSS DFF_X1 
Xprod_reg_27_ N27 n1_G3B1I3 p[27] SYNOPSYS_UNCONNECTED_85 VDD VSS DFF_X1 
Xprod_reg_28_ N28 n1_G3B1I3 p[28] SYNOPSYS_UNCONNECTED_84 VDD VSS DFF_X1 
Xprod_reg_29_ N29 n1_G3B1I4 p[29] SYNOPSYS_UNCONNECTED_83 VDD VSS DFF_X1 
Xprod_reg_30_ N30 n1 p[30] SYNOPSYS_UNCONNECTED_82 VDD VSS DFF_X1 
Xprod_reg_31_ N31 n1 p[31] SYNOPSYS_UNCONNECTED_81 VDD VSS DFF_X1 
Xprod_reg_32_ N32 clk p[32] SYNOPSYS_UNCONNECTED_80 VDD VSS DFF_X1 
Xb_reg_reg_0_ b[0] clk b_reg[0] SYNOPSYS_UNCONNECTED_79 VDD VSS DFF_X1 
Xb_reg_reg_1_ b[1] clk b_reg[1] SYNOPSYS_UNCONNECTED_78 VDD VSS DFF_X1 
Xb_reg_reg_2_ b[2] n2_G3B1I1 b_reg[2] SYNOPSYS_UNCONNECTED_77 VDD VSS DFF_X1 
Xb_reg_reg_3_ b[3] n2_G3B1I2 b_reg[3] SYNOPSYS_UNCONNECTED_76 VDD VSS DFF_X1 
Xb_reg_reg_4_ b[4] n2_G3B1I4 b_reg[4] SYNOPSYS_UNCONNECTED_75 VDD VSS DFF_X1 
Xb_reg_reg_5_ b[5] n1_G3B1I3 b_reg[5] SYNOPSYS_UNCONNECTED_74 VDD VSS DFF_X1 
Xb_reg_reg_6_ b[6] n1_G3B1I3 b_reg[6] SYNOPSYS_UNCONNECTED_73 VDD VSS DFF_X1 
Xb_reg_reg_7_ b[7] n1_G3B1I2 b_reg[7] SYNOPSYS_UNCONNECTED_72 VDD VSS DFF_X1 
Xb_reg_reg_8_ b[8] n1_G3B1I3 b_reg[8] SYNOPSYS_UNCONNECTED_71 VDD VSS DFF_X1 
Xb_reg_reg_9_ b[9] n1_G3B1I3 b_reg[9] SYNOPSYS_UNCONNECTED_70 VDD VSS DFF_X1 
Xb_reg_reg_10_ b[10] n1_G3B1I3 b_reg[10] SYNOPSYS_UNCONNECTED_69 VDD VSS DFF_X1 
Xb_reg_reg_11_ b[11] n1_G3B1I4 b_reg[11] SYNOPSYS_UNCONNECTED_68 VDD VSS DFF_X1 
Xb_reg_reg_12_ b[12] n1_G3B1I4 b_reg[12] SYNOPSYS_UNCONNECTED_67 VDD VSS DFF_X1 
Xb_reg_reg_13_ b[13] n1_G3B1I4 b_reg[13] SYNOPSYS_UNCONNECTED_66 VDD VSS DFF_X1 
Xb_reg_reg_14_ b[14] n1 b_reg[14] SYNOPSYS_UNCONNECTED_65 VDD VSS DFF_X1 
Xb_reg_reg_15_ b[15] n1 b_reg[15] SYNOPSYS_UNCONNECTED_64 VDD VSS DFF_X1 
Xb_reg_reg_16_ b[16] n1 b_reg[16] SYNOPSYS_UNCONNECTED_63 VDD VSS DFF_X1 
Xb_reg_reg_17_ b[17] n2_G3B1I4 b_reg[17] SYNOPSYS_UNCONNECTED_62 VDD VSS DFF_X1 
Xa_reg_reg_0_ a[0] n2_G3B1I2 a_reg[0] SYNOPSYS_UNCONNECTED_61 VDD VSS DFF_X1 
Xa_reg_reg_1_ a[1] n2_G3B1I1 a_reg[1] SYNOPSYS_UNCONNECTED_60 VDD VSS DFF_X1 
Xa_reg_reg_2_ a[2] n2_G3B1I2 a_reg[2] SYNOPSYS_UNCONNECTED_59 VDD VSS DFF_X1 
Xa_reg_reg_3_ a[3] n2_G3B1I2 a_reg[3] SYNOPSYS_UNCONNECTED_58 VDD VSS DFF_X1 
Xa_reg_reg_4_ a[4] n2_G3B1I2 a_reg[4] SYNOPSYS_UNCONNECTED_57 VDD VSS DFF_X1 
Xa_reg_reg_5_ a[5] n2_G3B1I1 a_reg[5] SYNOPSYS_UNCONNECTED_56 VDD VSS DFF_X1 
Xa_reg_reg_6_ a[6] n2_G3B1I4 a_reg[6] SYNOPSYS_UNCONNECTED_55 VDD VSS DFF_X1 
Xa_reg_reg_7_ a[7] n2_G3B1I4 a_reg[7] SYNOPSYS_UNCONNECTED_54 VDD VSS DFF_X1 
Xa_reg_reg_8_ a[8] n2_G3B1I4 a_reg[8] SYNOPSYS_UNCONNECTED_53 VDD VSS DFF_X1 
Xa_reg_reg_9_ a[9] n1 a_reg[9] SYNOPSYS_UNCONNECTED_52 VDD VSS DFF_X1 
Xa_reg_reg_10_ a[10] n2_G3B1I1 a_reg[10] SYNOPSYS_UNCONNECTED_51 VDD VSS DFF_X1 
Xa_reg_reg_11_ a[11] n2_G3B1I1 a_reg[11] SYNOPSYS_UNCONNECTED_50 VDD VSS DFF_X1 
Xa_reg_reg_12_ a[12] n2_G3B1I4 a_reg[12] SYNOPSYS_UNCONNECTED_49 VDD VSS DFF_X1 
Xa_reg_reg_13_ a[13] n2_G3B1I4 a_reg[13] SYNOPSYS_UNCONNECTED_48 VDD VSS DFF_X1 
Xa_reg_reg_14_ a[14] n2_G3B1I4 a_reg[14] SYNOPSYS_UNCONNECTED_47 VDD VSS DFF_X1 
Xa_reg_reg_15_ LOGIC0_X1_U0_net n2_G3B1I2 a_reg[15] SYNOPSYS_UNCONNECTED_46 VDD 
+ VSS DFF_X1 
XU1 clk n1 VDD VSS BUF_X32 
XCLKBUF_X1_G3B1I21 n1 n1_G3B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G3B1I4 clk n2_G3B1I4 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I31 n1 n1_G3B1I3 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I41 n1 n1_G3B1I4 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I1 clk n2_G3B1I1 VDD VSS CLKBUF_X2 
XCLKBUF_X1_G3B1I2 clk n2_G3B1I2 VDD VSS CLKBUF_X2 
Xmult_60 N33 N32 N31 N30 N29 N28 N27 N26 N25 N24 N23 N22 N21 N20 N19 N18 N17 N16 
+ N15 N14 N13 N12 N11 N101 N9 N8 N7 N6 N5 N4 N3 N2 N100 N0 VDD VDD VSS b_reg[17] 
+ b_reg[16] b_reg[15] b_reg[14] b_reg[13] b_reg[12] b_reg[11] b_reg[10] b_reg[9] 
+ b_reg[8] b_reg[7] b_reg[6] b_reg[5] b_reg[4] b_reg[3] b_reg[2] b_reg[1] b_reg[0] 
+ a_reg[15] a_reg[14] a_reg[13] a_reg[12] a_reg[11] a_reg[10] a_reg[9] a_reg[8] 
+ a_reg[7] a_reg[6] a_reg[5] a_reg[4] a_reg[3] a_reg[2] a_reg[1] a_reg[0] gng_smul_16_18_DW02_mult_0 
.ENDS

.SUBCKT gng_interp clk rstn valid_in valid_out VDD VSS IN0 IN1 data_out[15] data_out[14] 
+ data_out[13] data_out[12] data_out[11] data_out[10] data_out[9] data_out[8] data_out[7] 
+ data_out[6] data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] 
+ data_in[63] data_in[62] data_in[61] data_in[60] data_in[59] data_in[58] data_in[57] 
+ data_in[56] data_in[55] data_in[54] data_in[53] data_in[52] data_in[51] data_in[50] 
+ data_in[49] data_in[48] data_in[47] data_in[46] data_in[45] data_in[44] data_in[43] 
+ data_in[42] data_in[41] data_in[40] data_in[39] data_in[38] data_in[37] data_in[36] 
+ data_in[35] data_in[34] data_in[33] data_in[32] data_in[31] data_in[30] data_in[29] 
+ data_in[28] data_in[27] data_in[26] data_in[25] data_in[24] data_in[23] data_in[22] 
+ data_in[21] data_in[20] data_in[19] data_in[18] data_in[17] data_in[16] data_in[15] 
+ data_in[14] data_in[13] data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] 
+ data_in[7] data_in[6] data_in[5] data_in[4] data_in[3] data_in[2] data_in[1] data_in[0] 
+ IN2 clk_cts_3 
XU153 n132 n7310 VDD VSS CLKBUF_X2 
XU152 n204 n7210 VDD VSS BUF_X1 
XU150 n142 n7011 VDD VSS BUF_X2 
XU148 n208 n6810 VDD VSS BUF_X2 
Xx_r2_reg_7_ n1303 n10_G2B1I4 x_r2[7] SYNOPSYS_UNCONNECTED_539 VDD VSS DFF_X1 
Xx_r1_reg_7_ n201 n6_G2B1I4 x_r1[7] SYNOPSYS_UNCONNECTED_538 VDD VSS DFF_X1 
Xx_r3_reg_8_ n1293 n10_G2B1I3 x_r3[8] SYNOPSYS_UNCONNECTED_537 VDD VSS DFF_X1 
Xx_r2_reg_8_ n209 n10_G2B1I4 x_r2[8] SYNOPSYS_UNCONNECTED_536 VDD VSS DFF_X1 
Xx_r1_reg_8_ n1334 n60 x_r1[8] SYNOPSYS_UNCONNECTED_535 VDD VSS DFF_X1 
Xx_r3_reg_9_ n1280 n8_G2B1I2 x_r3[9] SYNOPSYS_UNCONNECTED_534 VDD VSS DFF_X1 
Xx_r2_reg_9_ n1276 n8_G2B1I7 x_r2[9] SYNOPSYS_UNCONNECTED_533 VDD VSS DFF_X1 
Xx_r1_reg_9_ n1307 n8_G2B1I2 x_r1[9] SYNOPSYS_UNCONNECTED_532 VDD VSS DFF_X1 
Xx_r3_reg_10_ n1266 n10_G2B1I4 x_r3[10] SYNOPSYS_UNCONNECTED_531 VDD VSS DFF_X1 
Xx_r2_reg_10_ n1262 n6_G2B1I5 x_r2[10] SYNOPSYS_UNCONNECTED_530 VDD VSS DFF_X1 
Xx_r1_reg_10_ n200 n6_G2B1I4 x_r1[10] SYNOPSYS_UNCONNECTED_529 VDD VSS DFF_X1 
Xx_r3_reg_11_ n1253 n10_G2B1I4 x_r3[11] SYNOPSYS_UNCONNECTED_528 VDD VSS DFF_X1 
Xx_r2_reg_11_ n1249 n6_G2B1I5 x_r2[11] SYNOPSYS_UNCONNECTED_527 VDD VSS DFF_X1 
Xx_r1_reg_11_ n198 n6_G2B1I4 x_r1[11] SYNOPSYS_UNCONNECTED_526 VDD VSS DFF_X1 
Xx_r3_reg_12_ n1239 n10_G2B1I2 x_r3[12] SYNOPSYS_UNCONNECTED_525 VDD VSS DFF_X1 
Xx_r2_reg_12_ n1235 n10_G2B1I4 x_r2[12] SYNOPSYS_UNCONNECTED_524 VDD VSS DFF_X1 
Xx_r1_reg_12_ n1970 n6_G2B1I4 x_r1[12] SYNOPSYS_UNCONNECTED_523 VDD VSS DFF_X1 
Xx_r3_reg_13_ n1226 n10_G2B1I3 x_r3[13] SYNOPSYS_UNCONNECTED_522 VDD VSS DFF_X1 
Xx_r2_reg_13_ n1222 n10_G2B1I2 x_r2[13] SYNOPSYS_UNCONNECTED_521 VDD VSS DFF_X1 
Xx_r1_reg_13_ n1950 n6_G2B1I3 x_r1[13] SYNOPSYS_UNCONNECTED_520 VDD VSS DFF_X1 
Xx_r3_reg_14_ n1212 n10_G2B1I2 x_r3[14] SYNOPSYS_UNCONNECTED_519 VDD VSS DFF_X1 
Xx_r2_reg_14_ n1208 n10_G2B1I2 x_r2[14] SYNOPSYS_UNCONNECTED_518 VDD VSS DFF_X1 
Xx_r1_reg_14_ n1940 n6_G2B1I3 x_r1[14] SYNOPSYS_UNCONNECTED_517 VDD VSS DFF_X1 
Xx_reg_0_ n1195 n11_G2B1I7 SYNOPSYS_UNCONNECTED_516 n59 VDD VSS DFF_X1 
Xx_reg_1_ n1191 n11_G2B1I7 SYNOPSYS_UNCONNECTED_515 n6110 VDD VSS DFF_X1 
Xx_reg_2_ n1190 n11_G2B1I6 SYNOPSYS_UNCONNECTED_514 n630 VDD VSS DFF_X1 
Xx_reg_3_ N80 n11_G2B1I6 SYNOPSYS_UNCONNECTED_513 n650 VDD VSS DFF_X1 
Xx_reg_4_ n1186 n11_G2B1I1 SYNOPSYS_UNCONNECTED_512 n670 VDD VSS DFF_X1 
Xx_reg_5_ n1182 n11_G2B1I4 SYNOPSYS_UNCONNECTED_511 n690 VDD VSS DFF_X1 
Xx_reg_6_ n1178 n11_G2B1I5 SYNOPSYS_UNCONNECTED_510 n711 VDD VSS DFF_X1 
Xx_reg_7_ n1174 n11_G2B1I3 SYNOPSYS_UNCONNECTED_509 n730 VDD VSS DFF_X1 
Xx_reg_8_ n1167 n11_G2B1I6 SYNOPSYS_UNCONNECTED_508 n750 VDD VSS DFF_X1 
Xx_reg_9_ n1166 n2 SYNOPSYS_UNCONNECTED_507 n770 VDD VSS DFF_X1 
Xx_reg_10_ n1163 n11_G2B1I2 SYNOPSYS_UNCONNECTED_506 n790 VDD VSS DFF_X1 
Xx_reg_11_ n1159 n11_G2B1I3 SYNOPSYS_UNCONNECTED_505 n811 VDD VSS DFF_X1 
Xx_reg_12_ n1157 n11_G2B1I3 SYNOPSYS_UNCONNECTED_504 n830 VDD VSS DFF_X1 
Xx_reg_13_ n1153 n11_G2B1I3 SYNOPSYS_UNCONNECTED_503 n850 VDD VSS DFF_X1 
Xx_reg_14_ n1149 n11_G2B1I3 SYNOPSYS_UNCONNECTED_502 n870 VDD VSS DFF_X1 
Xoffset_reg_0_ n1142 n6 offset[0] SYNOPSYS_UNCONNECTED_501 VDD VSS DFF_X1 
Xoffset_reg_1_ n1141 n8_G2B1I7 offset[1] SYNOPSYS_UNCONNECTED_500 VDD VSS DFF_X1 
Xmask_reg_0_ n1134 n11_G2B1I7 SYNOPSYS_UNCONNECTED_499 n6000 VDD VSS DFF_X1 
Xmask_reg_1_ n1129 n11_G2B1I7 SYNOPSYS_UNCONNECTED_498 n6200 VDD VSS DFF_X1 
Xmask_reg_2_ N620 n11_G2B1I5 SYNOPSYS_UNCONNECTED_497 n640 VDD VSS DFF_X1 
Xmask_reg_3_ N63 n11_G2B1I6 SYNOPSYS_UNCONNECTED_496 n660 VDD VSS DFF_X1 
Xmask_reg_4_ n1109 n11_G2B1I6 SYNOPSYS_UNCONNECTED_495 n680 VDD VSS DFF_X1 
Xmask_reg_5_ n1103 n11_G2B1I5 SYNOPSYS_UNCONNECTED_494 n7000 VDD VSS DFF_X1 
Xmask_reg_6_ N66 n11_G2B1I5 SYNOPSYS_UNCONNECTED_493 n720 VDD VSS DFF_X1 
Xmask_reg_7_ N67 n11_G2B1I2 SYNOPSYS_UNCONNECTED_492 n740 VDD VSS DFF_X1 
Xmask_reg_8_ N68 n11_G2B1I6 SYNOPSYS_UNCONNECTED_491 n760 VDD VSS DFF_X1 
Xmask_reg_9_ N69 n11_G2B1I4 SYNOPSYS_UNCONNECTED_490 n780 VDD VSS DFF_X1 
Xmask_reg_10_ n1085 n6_G2B1I3 SYNOPSYS_UNCONNECTED_489 n800 VDD VSS DFF_X1 
Xmask_reg_11_ N71 n11_G2B1I2 SYNOPSYS_UNCONNECTED_488 n820 VDD VSS DFF_X1 
Xmask_reg_12_ N72 n11_G2B1I5 SYNOPSYS_UNCONNECTED_487 n840 VDD VSS DFF_X1 
Xmask_reg_13_ N73 n11_G2B1I2 SYNOPSYS_UNCONNECTED_486 n860 VDD VSS DFF_X1 
Xmask_reg_14_ n1083 n11_G2B1I2 SYNOPSYS_UNCONNECTED_485 n880 VDD VSS DFF_X1 
Xnum_lzd_r_reg_0_ n1920 n11_G2B1I4 num_lzd_r[0] n1110 VDD VSS DFF_X2 
Xnum_lzd_r_reg_1_ n1082 n11_G2B1I4 num_lzd_r[1] n1010 VDD VSS DFF_X1 
Xnum_lzd_r_reg_2_ n1081 n11_G2B1I4 num_lzd_r[2] n910 VDD VSS DFF_X1 
Xnum_lzd_r_reg_3_ n1079 n11_G2B1I3 num_lzd_r[3] n810 VDD VSS DFF_X1 
Xnum_lzd_r_reg_4_ n1075 n11_G2B1I4 num_lzd_r[4] n710 VDD VSS DFF_X1 
Xnum_lzd_r_reg_5_ n1073 n11_G2B1I4 num_lzd_r[5] SYNOPSYS_UNCONNECTED_484 VDD VSS DFF_X1 
Xc0_r2_reg_8_ n1071 n7_G2B1I1 c0_r2[8] SYNOPSYS_UNCONNECTED_483 VDD VSS DFF_X1 
Xc0_r1_reg_8_ c0[8] n7_G2B1I1 c0_r1[8] SYNOPSYS_UNCONNECTED_482 VDD VSS DFF_X1 
Xc0_r4_reg_9_ n1066 n7_G2B1I4 c0_r4[9] SYNOPSYS_UNCONNECTED_481 VDD VSS DFF_X1 
Xc0_r3_reg_9_ n1062 n7_G2B1I4 c0_r3[9] SYNOPSYS_UNCONNECTED_480 VDD VSS DFF_X1 
Xc0_r2_reg_9_ n1880 n7_G2B1I4 c0_r2[9] SYNOPSYS_UNCONNECTED_479 VDD VSS DFF_X1 
Xc0_r1_reg_9_ c0[9] n62 c0_r1[9] SYNOPSYS_UNCONNECTED_478 VDD VSS DFF_X1 
Xc0_r4_reg_10_ n1049 n62 c0_r4[10] SYNOPSYS_UNCONNECTED_477 VDD VSS DFF_X1 
Xc0_r3_reg_10_ n1048 n62_G2B1I2 c0_r3[10] SYNOPSYS_UNCONNECTED_476 VDD VSS DFF_X1 
Xc0_r2_reg_10_ n1044 n62_G2B1I2 c0_r2[10] SYNOPSYS_UNCONNECTED_475 VDD VSS DFF_X1 
Xc0_r1_reg_10_ c0[10] n63_G2B1I2 c0_r1[10] SYNOPSYS_UNCONNECTED_474 VDD VSS DFF_X1 
Xc0_r4_reg_11_ n1039 n6_G2B1I5 c0_r4[11] SYNOPSYS_UNCONNECTED_473 VDD VSS DFF_X1 
Xc0_r3_reg_11_ n1035 n6_G2B1I5 c0_r3[11] SYNOPSYS_UNCONNECTED_472 VDD VSS DFF_X1 
Xc0_r2_reg_11_ n1031 n6_G2B1I3 c0_r2[11] SYNOPSYS_UNCONNECTED_471 VDD VSS DFF_X1 
Xc0_r1_reg_11_ c0[11] n6_G2B1I3 c0_r1[11] SYNOPSYS_UNCONNECTED_470 VDD VSS DFF_X1 
Xc0_r4_reg_12_ n1026 n6_G2B1I5 c0_r4[12] SYNOPSYS_UNCONNECTED_469 VDD VSS DFF_X1 
Xc0_r3_reg_12_ n1022 n6_G2B1I3 c0_r3[12] SYNOPSYS_UNCONNECTED_468 VDD VSS DFF_X1 
Xc0_r2_reg_12_ n1870 n6_G2B1I3 c0_r2[12] SYNOPSYS_UNCONNECTED_467 VDD VSS DFF_X1 
Xc0_r1_reg_12_ c0[12] n6 c0_r1[12] SYNOPSYS_UNCONNECTED_466 VDD VSS DFF_X1 
Xc0_r4_reg_13_ n1013 n60_G2B1I5 c0_r4[13] SYNOPSYS_UNCONNECTED_465 VDD VSS DFF_X1 
Xc0_r3_reg_13_ n1007 n60_G2B1I5 c0_r3[13] SYNOPSYS_UNCONNECTED_464 VDD VSS DFF_X1 
Xc0_r2_reg_13_ n1003 n60_G2B1I5 c0_r2[13] SYNOPSYS_UNCONNECTED_463 VDD VSS DFF_X1 
Xc0_r1_reg_13_ c0[13] n11_G2B1I6 c0_r1[13] SYNOPSYS_UNCONNECTED_462 VDD VSS DFF_X1 
Xc0_r4_reg_14_ n998 n8_G2B1I2 c0_r4[14] SYNOPSYS_UNCONNECTED_461 VDD VSS DFF_X1 
Xc0_r3_reg_14_ n994 n8_G2B1I7 c0_r3[14] SYNOPSYS_UNCONNECTED_460 VDD VSS DFF_X1 
Xc0_r2_reg_14_ n989 n8_G2B1I7 c0_r2[14] SYNOPSYS_UNCONNECTED_459 VDD VSS DFF_X1 
Xc0_r1_reg_14_ c0[14] n8_G2B1I7 c0_r1[14] SYNOPSYS_UNCONNECTED_458 VDD VSS DFF_X1 
Xc0_r4_reg_15_ n985 n11_G2B1I1 c0_r4[15] SYNOPSYS_UNCONNECTED_457 VDD VSS DFF_X1 
Xc0_r3_reg_15_ n981 n60_G2B1I1 c0_r3[15] SYNOPSYS_UNCONNECTED_456 VDD VSS DFF_X1 
Xc0_r2_reg_15_ n976 n60_G2B1I1 c0_r2[15] SYNOPSYS_UNCONNECTED_455 VDD VSS DFF_X1 
Xc0_r1_reg_15_ c0[15] n60_G2B1I5 c0_r1[15] SYNOPSYS_UNCONNECTED_454 VDD VSS DFF_X1 
Xc0_r4_reg_16_ n972 n8_G2B1I7 c0_r4[16] SYNOPSYS_UNCONNECTED_453 VDD VSS DFF_X1 
Xc0_r3_reg_16_ n968 n8_G2B1I1 c0_r3[16] SYNOPSYS_UNCONNECTED_452 VDD VSS DFF_X1 
Xc0_r2_reg_16_ n964 n8_G2B1I1 c0_r2[16] SYNOPSYS_UNCONNECTED_451 VDD VSS DFF_X1 
Xc0_r1_reg_16_ c0[16] n8_G2B1I1 c0_r1[16] SYNOPSYS_UNCONNECTED_450 VDD VSS DFF_X1 
Xc0_r4_reg_17_ n960 n11_G2B1I1 c0_r4[17] SYNOPSYS_UNCONNECTED_449 VDD VSS DFF_X1 
Xc0_r3_reg_17_ n956 n11_G2B1I1 c0_r3[17] SYNOPSYS_UNCONNECTED_448 VDD VSS DFF_X1 
Xc0_r2_reg_17_ n952 n11_G2B1I1 c0_r2[17] SYNOPSYS_UNCONNECTED_447 VDD VSS DFF_X1 
Xc0_r1_reg_17_ c0[17] n11_G2B1I6 c0_r1[17] SYNOPSYS_UNCONNECTED_446 VDD VSS DFF_X1 
Xc1_r1_reg_0_ c1[0] n11_G2B1I5 c1_r1[0] SYNOPSYS_UNCONNECTED_445 VDD VSS DFF_X1 
Xc1_r1_reg_1_ c1[1] n6_G2B1I3 c1_r1[1] SYNOPSYS_UNCONNECTED_444 VDD VSS DFF_X1 
Xc1_r1_reg_2_ c1[2] n6 c1_r1[2] SYNOPSYS_UNCONNECTED_443 VDD VSS DFF_X1 
Xc1_r1_reg_3_ c1[3] n6_G2B1I3 c1_r1[3] SYNOPSYS_UNCONNECTED_442 VDD VSS DFF_X1 
Xc1_r1_reg_4_ c1[4] n6_G2B1I5 c1_r1[4] SYNOPSYS_UNCONNECTED_441 VDD VSS DFF_X1 
Xc1_r1_reg_5_ c1[5] n62_G2B1I2 c1_r1[5] SYNOPSYS_UNCONNECTED_440 VDD VSS DFF_X1 
Xc1_r1_reg_6_ c1[6] n62_G2B1I2 c1_r1[6] SYNOPSYS_UNCONNECTED_439 VDD VSS DFF_X1 
Xc1_r1_reg_7_ c1[7] n62 c1_r1[7] SYNOPSYS_UNCONNECTED_438 VDD VSS DFF_X1 
Xc1_r1_reg_8_ c1[8] n7_G2B1I4 c1_r1[8] SYNOPSYS_UNCONNECTED_437 VDD VSS DFF_X1 
Xc1_r1_reg_9_ c1[9] n7_G2B1I4 c1_r1[9] SYNOPSYS_UNCONNECTED_436 VDD VSS DFF_X1 
Xc1_r1_reg_10_ c1[10] n7_G2B1I4 c1_r1[10] SYNOPSYS_UNCONNECTED_435 VDD VSS DFF_X1 
Xc1_r1_reg_11_ c1[11] n62 c1_r1[11] SYNOPSYS_UNCONNECTED_434 VDD VSS DFF_X1 
Xc1_r1_reg_12_ c1[12] n62_G2B1I2 c1_r1[12] SYNOPSYS_UNCONNECTED_433 VDD VSS DFF_X1 
Xc1_r1_reg_13_ c1[13] n62_G2B1I2 c1_r1[13] SYNOPSYS_UNCONNECTED_432 VDD VSS DFF_X1 
Xc1_r1_reg_14_ c1[14] n63_G2B1I8 c1_r1[14] SYNOPSYS_UNCONNECTED_431 VDD VSS DFF_X1 
Xc1_r1_reg_15_ c1[15] n63_G2B1I8 c1_r1[15] SYNOPSYS_UNCONNECTED_430 VDD VSS DFF_X1 
Xc1_r1_reg_16_ c1[16] n63_G2B1I8 c1_r1[16] SYNOPSYS_UNCONNECTED_429 VDD VSS DFF_X1 
Xc1_r1_reg_17_ c1[17] n63_G2B1I8 c1_r1[17] SYNOPSYS_UNCONNECTED_428 VDD VSS DFF_X1 
Xx_r4_reg_0_ n947 n6_G2B1I2 x_r4[0] SYNOPSYS_UNCONNECTED_427 VDD VSS DFF_X1 
Xx_r4_reg_1_ n943 n6_G2B1I2 x_r4[1] SYNOPSYS_UNCONNECTED_426 VDD VSS DFF_X1 
Xx_r4_reg_2_ n938 n10_G2B1I3 x_r4[2] SYNOPSYS_UNCONNECTED_425 VDD VSS DFF_X1 
Xx_r4_reg_3_ n934 n6_G2B1I2 x_r4[3] SYNOPSYS_UNCONNECTED_424 VDD VSS DFF_X1 
Xx_r4_reg_4_ n1860 n61_G2B1I1 x_r4[4] SYNOPSYS_UNCONNECTED_423 VDD VSS DFF_X1 
Xx_r4_reg_5_ n925 n6_G2B1I2 x_r4[5] SYNOPSYS_UNCONNECTED_422 VDD VSS DFF_X1 
Xx_r4_reg_6_ n1850 n61_G2B1I1 x_r4[6] SYNOPSYS_UNCONNECTED_421 VDD VSS DFF_X1 
Xx_r4_reg_7_ n916 n61_G2B1I1 x_r4[7] SYNOPSYS_UNCONNECTED_420 VDD VSS DFF_X1 
Xx_r4_reg_8_ n912 n61_G2B1I1 x_r4[8] SYNOPSYS_UNCONNECTED_419 VDD VSS DFF_X1 
Xx_r4_reg_9_ n906 n8_G2B1I2 x_r4[9] SYNOPSYS_UNCONNECTED_418 VDD VSS DFF_X1 
Xx_r4_reg_10_ n902 n10_G2B1I2 x_r4[10] SYNOPSYS_UNCONNECTED_417 VDD VSS DFF_X1 
Xx_r4_reg_11_ n897 n10_G2B1I2 x_r4[11] SYNOPSYS_UNCONNECTED_416 VDD VSS DFF_X1 
Xx_r4_reg_12_ n893 n10_G2B1I3 x_r4[12] SYNOPSYS_UNCONNECTED_415 VDD VSS DFF_X1 
Xx_r4_reg_13_ n888 n10_G2B1I3 x_r4[13] SYNOPSYS_UNCONNECTED_414 VDD VSS DFF_X1 
Xx_r4_reg_14_ n884 n10_G2B1I3 x_r4[14] SYNOPSYS_UNCONNECTED_413 VDD VSS DFF_X1 
Xx_r3_reg_0_ n879 n6_G2B1I2 x_r3[0] SYNOPSYS_UNCONNECTED_412 VDD VSS DFF_X1 
Xx_r2_reg_0_ n875 n6_G2B1I4 x_r2[0] SYNOPSYS_UNCONNECTED_411 VDD VSS DFF_X1 
Xx_r1_reg_0_ n141 n11_G2B1I5 x_r1[0] SYNOPSYS_UNCONNECTED_410 VDD VSS DFF_X1 
Xx_r3_reg_1_ n864 n6_G2B1I4 x_r3[1] SYNOPSYS_UNCONNECTED_409 VDD VSS DFF_X1 
Xx_r2_reg_1_ n859 n6_G2B1I4 x_r2[1] SYNOPSYS_UNCONNECTED_408 VDD VSS DFF_X1 
Xx_r1_reg_1_ n1840 n11_G2B1I6 x_r1[1] SYNOPSYS_UNCONNECTED_407 VDD VSS DFF_X1 
Xx_r3_reg_2_ n849 n10_G2B1I4 x_r3[2] SYNOPSYS_UNCONNECTED_406 VDD VSS DFF_X1 
Xx_r2_reg_2_ n845 n6_G2B1I2 x_r2[2] SYNOPSYS_UNCONNECTED_405 VDD VSS DFF_X1 
Xx_r1_reg_2_ n1820 n6_G2B1I4 x_r1[2] SYNOPSYS_UNCONNECTED_404 VDD VSS DFF_X1 
Xx_r3_reg_3_ n181 n6_G2B1I4 x_r3[3] SYNOPSYS_UNCONNECTED_403 VDD VSS DFF_X1 
Xx_r2_reg_3_ n829 n60 x_r2[3] SYNOPSYS_UNCONNECTED_402 VDD VSS DFF_X1 
Xx_r1_reg_3_ n180 n60_G2B1I5 x_r1[3] SYNOPSYS_UNCONNECTED_401 VDD VSS DFF_X1 
Xx_r3_reg_4_ n819 n10_G2B1I1 x_r3[4] SYNOPSYS_UNCONNECTED_400 VDD VSS DFF_X1 
Xx_r2_reg_4_ n815 n6_G2B1I2 x_r2[4] SYNOPSYS_UNCONNECTED_399 VDD VSS DFF_X1 
Xx_r1_reg_4_ n178 n60_G2B1I5 x_r1[4] SYNOPSYS_UNCONNECTED_398 VDD VSS DFF_X1 
Xx_r3_reg_5_ n804 n6_G2B1I2 x_r3[5] SYNOPSYS_UNCONNECTED_397 VDD VSS DFF_X1 
Xx_r2_reg_5_ n210 n6_G2B1I2 x_r2[5] SYNOPSYS_UNCONNECTED_396 VDD VSS DFF_X1 
Xx_r1_reg_5_ n176 n60 x_r1[5] SYNOPSYS_UNCONNECTED_395 VDD VSS DFF_X1 
Xx_r3_reg_6_ n789 n10_G2B1I1 x_r3[6] SYNOPSYS_UNCONNECTED_394 VDD VSS DFF_X1 
Xx_r2_reg_6_ n785 n10_G2B1I4 x_r2[6] SYNOPSYS_UNCONNECTED_393 VDD VSS DFF_X1 
Xx_r1_reg_6_ n175 n6_G2B1I4 x_r1[6] SYNOPSYS_UNCONNECTED_392 VDD VSS DFF_X1 
Xx_r3_reg_7_ n775 n10_G2B1I3 x_r3[7] SYNOPSYS_UNCONNECTED_391 VDD VSS DFF_X1 
Xsum2_rnd_reg_8_ n173 n62_G2B1I2 SYNOPSYS_UNCONNECTED_390 n35 VDD VSS DFF_X1 
Xsum2_rnd_reg_9_ n171 n62_G2B1I2 SYNOPSYS_UNCONNECTED_389 n34 VDD VSS DFF_X1 
Xsum2_rnd_reg_10_ n755 n60 SYNOPSYS_UNCONNECTED_388 n33 VDD VSS DFF_X1 
Xsum2_rnd_reg_11_ n170 n60_G2B1I1 SYNOPSYS_UNCONNECTED_387 n32 VDD VSS DFF_X1 
Xsum2_rnd_reg_12_ n169 n60_G2B1I1 SYNOPSYS_UNCONNECTED_386 n31 VDD VSS DFF_X1 
Xsum2_rnd_reg_13_ n168 n11_G2B1I7 SYNOPSYS_UNCONNECTED_385 n30 VDD VSS DFF_X1 
Xsum2_rnd_reg_14_ n167 n2 SYNOPSYS_UNCONNECTED_384 n29 VDD VSS DFF_X1 
Xsum2_reg_2_ N116 n7 sum2[2] SYNOPSYS_UNCONNECTED_383 VDD VSS DFF_X1 
Xsum2_reg_3_ N117 n7 sum2[3] SYNOPSYS_UNCONNECTED_382 VDD VSS DFF_X1 
Xsum2_reg_4_ N118 n9_G2B1I2 sum2[4] SYNOPSYS_UNCONNECTED_381 VDD VSS DFF_X1 
Xsum2_reg_5_ N119 n9_G2B1I2 sum2[5] SYNOPSYS_UNCONNECTED_380 VDD VSS DFF_X1 
Xsum2_reg_6_ N120 n9_G2B1I2 sum2[6] SYNOPSYS_UNCONNECTED_379 VDD VSS DFF_X1 
Xsum2_reg_7_ n1336 n7_G2B1I2 sum2[7] SYNOPSYS_UNCONNECTED_378 VDD VSS DFF_X1 
Xsum2_reg_8_ N122 n7 sum2[8] SYNOPSYS_UNCONNECTED_377 VDD VSS DFF_X1 
Xsum2_reg_9_ N123 n7 sum2[9] SYNOPSYS_UNCONNECTED_376 VDD VSS DFF_X1 
Xsum2_reg_10_ N124 n62 sum2[10] SYNOPSYS_UNCONNECTED_375 VDD VSS DFF_X1 
Xsum2_reg_11_ N125 n62_G2B1I2 sum2[11] SYNOPSYS_UNCONNECTED_374 VDD VSS DFF_X1 
Xsum2_reg_12_ N126 n63_G2B1I2 sum2[12] SYNOPSYS_UNCONNECTED_373 VDD VSS DFF_X1 
Xsum2_reg_13_ n1305 n60_G2B1I5 sum2[13] SYNOPSYS_UNCONNECTED_372 VDD VSS DFF_X1 
Xsum2_reg_14_ N128 n60_G2B1I1 sum2[14] SYNOPSYS_UNCONNECTED_371 VDD VSS DFF_X1 
Xsum2_reg_15_ N129 n60_G2B1I1 sum2[15] SYNOPSYS_UNCONNECTED_370 VDD VSS DFF_X1 
Xsum2_reg_16_ N130 n11_G2B1I7 sum2[16] SYNOPSYS_UNCONNECTED_369 VDD VSS DFF_X1 
Xsum2_reg_17_ N131 n11_G2B1I7 SYNOPSYS_UNCONNECTED_368 n58 VDD VSS DFF_X1 
Xvalid_in_r_reg_8_ n732 n8_G2B1I4 valid_in_r[8] SYNOPSYS_UNCONNECTED_367 VDD VSS DFF_X1 
Xvalid_in_r_reg_7_ n727 n8_G2B1I5 valid_in_r[7] SYNOPSYS_UNCONNECTED_366 VDD VSS DFF_X1 
Xvalid_in_r_reg_6_ n723 n8_G2B1I8 valid_in_r[6] SYNOPSYS_UNCONNECTED_365 VDD VSS DFF_X1 
Xvalid_in_r_reg_5_ n718 n8_G2B1I8 valid_in_r[5] SYNOPSYS_UNCONNECTED_364 VDD VSS DFF_X1 
Xvalid_in_r_reg_4_ n714 n8_G2B1I1 valid_in_r[4] SYNOPSYS_UNCONNECTED_363 VDD VSS DFF_X1 
Xvalid_in_r_reg_3_ n708 n8_G2B1I1 valid_in_r[3] SYNOPSYS_UNCONNECTED_362 VDD VSS DFF_X1 
Xvalid_in_r_reg_2_ N109 n8_G2B1I7 valid_in_r[2] SYNOPSYS_UNCONNECTED_361 VDD VSS DFF_X1 
Xvalid_in_r_reg_1_ n699 n2 valid_in_r[1] SYNOPSYS_UNCONNECTED_360 VDD VSS DFF_X1 
Xvalid_in_r_reg_0_ n692 n2 valid_in_r[0] SYNOPSYS_UNCONNECTED_359 VDD VSS DFF_X1 
Xsign_r_reg_8_ n691 n2 sign_r[8] n12 VDD VSS DFF_X1 
Xsign_r_reg_7_ n686 n2 sign_r[7] SYNOPSYS_UNCONNECTED_358 VDD VSS DFF_X1 
Xsign_r_reg_6_ n678 n2 sign_r[6] SYNOPSYS_UNCONNECTED_357 VDD VSS DFF_X1 
Xsign_r_reg_5_ n677 n2_G2B1I3 sign_r[5] SYNOPSYS_UNCONNECTED_356 VDD VSS DFF_X1 
Xsign_r_reg_4_ n673 n2_G2B1I3 sign_r[4] SYNOPSYS_UNCONNECTED_355 VDD VSS DFF_X1 
Xsign_r_reg_3_ n668 n2_G2B1I3 sign_r[3] SYNOPSYS_UNCONNECTED_354 VDD VSS DFF_X1 
Xsign_r_reg_2_ n664 n2_G2B1I3 sign_r[2] SYNOPSYS_UNCONNECTED_353 VDD VSS DFF_X1 
Xsign_r_reg_1_ n659 n2_G2B1I3 sign_r[1] SYNOPSYS_UNCONNECTED_352 VDD VSS DFF_X1 
Xsign_r_reg_0_ data_in[0] n2_G2B1I3 sign_r[0] SYNOPSYS_UNCONNECTED_351 VDD VSS DFF_X1 
Xc0_r5_reg_0_ n655 n8_G2B1I5 c0_r5[0] SYNOPSYS_UNCONNECTED_350 VDD VSS DFF_X1 
Xc0_r5_reg_1_ n651 n8_G2B1I5 c0_r5[1] SYNOPSYS_UNCONNECTED_349 VDD VSS DFF_X1 
Xc0_r5_reg_2_ n646 n8_G2B1I6 c0_r5[2] SYNOPSYS_UNCONNECTED_348 VDD VSS DFF_X1 
Xc0_r5_reg_3_ n642 n8_G2B1I6 c0_r5[3] SYNOPSYS_UNCONNECTED_347 VDD VSS DFF_X1 
Xc0_r5_reg_4_ n637 n7_G2B1I2 c0_r5[4] SYNOPSYS_UNCONNECTED_346 VDD VSS DFF_X1 
Xc0_r5_reg_5_ n633 n9_G2B1I2 c0_r5[5] SYNOPSYS_UNCONNECTED_345 VDD VSS DFF_X1 
Xc0_r5_reg_6_ n628 n9_G2B1I1 c0_r5[6] SYNOPSYS_UNCONNECTED_344 VDD VSS DFF_X1 
Xc0_r5_reg_7_ n624 n7_G2B1I1 c0_r5[7] SYNOPSYS_UNCONNECTED_343 VDD VSS DFF_X1 
Xc0_r5_reg_8_ n619 n7_G2B1I4 c0_r5[8] SYNOPSYS_UNCONNECTED_342 VDD VSS DFF_X1 
Xc0_r5_reg_9_ n615 n7_G2B1I4 c0_r5[9] SYNOPSYS_UNCONNECTED_341 VDD VSS DFF_X1 
Xc0_r5_reg_10_ n609 n62 c0_r5[10] SYNOPSYS_UNCONNECTED_340 VDD VSS DFF_X1 
Xc0_r5_reg_11_ n605 n6_G2B1I5 c0_r5[11] SYNOPSYS_UNCONNECTED_339 VDD VSS DFF_X1 
Xc0_r5_reg_12_ n601 n6_G2B1I5 c0_r5[12] SYNOPSYS_UNCONNECTED_338 VDD VSS DFF_X1 
Xc0_r5_reg_13_ n596 n60_G2B1I5 c0_r5[13] SYNOPSYS_UNCONNECTED_337 VDD VSS DFF_X1 
Xc0_r5_reg_14_ n140 n2 c0_r5[14] SYNOPSYS_UNCONNECTED_336 VDD VSS DFF_X1 
Xc0_r5_reg_15_ n588 n11_G2B1I1 c0_r5[15] SYNOPSYS_UNCONNECTED_335 VDD VSS DFF_X1 
Xc0_r5_reg_16_ n584 n8_G2B1I7 c0_r5[16] SYNOPSYS_UNCONNECTED_334 VDD VSS DFF_X1 
Xc0_r5_reg_17_ n580 n11_G2B1I1 c0_r5[17] SYNOPSYS_UNCONNECTED_333 VDD VSS DFF_X1 
Xc0_r4_reg_0_ n576 n8_G2B1I5 c0_r4[0] SYNOPSYS_UNCONNECTED_332 VDD VSS DFF_X1 
Xc0_r3_reg_0_ n572 n8_G2B1I5 c0_r3[0] SYNOPSYS_UNCONNECTED_331 VDD VSS DFF_X1 
Xc0_r2_reg_0_ n568 n8_G2B1I8 c0_r2[0] SYNOPSYS_UNCONNECTED_330 VDD VSS DFF_X1 
Xc0_r1_reg_0_ c0[0] n8_G2B1I8 c0_r1[0] SYNOPSYS_UNCONNECTED_329 VDD VSS DFF_X1 
Xc0_r4_reg_1_ n564 n8_G2B1I5 c0_r4[1] SYNOPSYS_UNCONNECTED_328 VDD VSS DFF_X1 
Xc0_r3_reg_1_ n560 n8_G2B1I8 c0_r3[1] SYNOPSYS_UNCONNECTED_327 VDD VSS DFF_X1 
Xc0_r2_reg_1_ n556 n8_G2B1I8 c0_r2[1] SYNOPSYS_UNCONNECTED_326 VDD VSS DFF_X1 
Xc0_r1_reg_1_ c0[1] n8_G2B1I8 c0_r1[1] SYNOPSYS_UNCONNECTED_325 VDD VSS DFF_X1 
Xc0_r4_reg_2_ n552 n8_G2B1I6 c0_r4[2] SYNOPSYS_UNCONNECTED_324 VDD VSS DFF_X1 
Xc0_r3_reg_2_ n548 n8_G2B1I6 c0_r3[2] SYNOPSYS_UNCONNECTED_323 VDD VSS DFF_X1 
Xc0_r2_reg_2_ n544 n8_G2B1I4 c0_r2[2] SYNOPSYS_UNCONNECTED_322 VDD VSS DFF_X1 
Xc0_r1_reg_2_ c0[2] n8_G2B1I4 c0_r1[2] SYNOPSYS_UNCONNECTED_321 VDD VSS DFF_X1 
Xc0_r4_reg_3_ n540 n8_G2B1I6 c0_r4[3] SYNOPSYS_UNCONNECTED_320 VDD VSS DFF_X1 
Xc0_r3_reg_3_ n536 n8_G2B1I4 c0_r3[3] SYNOPSYS_UNCONNECTED_319 VDD VSS DFF_X1 
Xc0_r2_reg_3_ n532 n8_G2B1I4 c0_r2[3] SYNOPSYS_UNCONNECTED_318 VDD VSS DFF_X1 
Xc0_r1_reg_3_ c0[3] n8_G2B1I4 c0_r1[3] SYNOPSYS_UNCONNECTED_317 VDD VSS DFF_X1 
Xc0_r4_reg_4_ n528 n7_G2B1I2 c0_r4[4] SYNOPSYS_UNCONNECTED_316 VDD VSS DFF_X1 
Xc0_r3_reg_4_ n524 n7_G2B1I2 c0_r3[4] SYNOPSYS_UNCONNECTED_315 VDD VSS DFF_X1 
Xc0_r2_reg_4_ n520 n7_G2B1I1 c0_r2[4] SYNOPSYS_UNCONNECTED_314 VDD VSS DFF_X1 
Xc0_r1_reg_4_ c0[4] n7_G2B1I1 c0_r1[4] SYNOPSYS_UNCONNECTED_313 VDD VSS DFF_X1 
Xc0_r4_reg_5_ n516 n9_G2B1I2 c0_r4[5] SYNOPSYS_UNCONNECTED_312 VDD VSS DFF_X1 
Xc0_r3_reg_5_ n512 n9_G2B1I2 c0_r3[5] SYNOPSYS_UNCONNECTED_311 VDD VSS DFF_X1 
Xc0_r2_reg_5_ n508 n7_G2B1I2 c0_r2[5] SYNOPSYS_UNCONNECTED_310 VDD VSS DFF_X1 
Xc0_r1_reg_5_ c0[5] n7_G2B1I1 c0_r1[5] SYNOPSYS_UNCONNECTED_309 VDD VSS DFF_X1 
Xc0_r4_reg_6_ n504 n9_G2B1I1 c0_r4[6] SYNOPSYS_UNCONNECTED_308 VDD VSS DFF_X1 
Xc0_r3_reg_6_ n500 n9_G2B1I1 c0_r3[6] SYNOPSYS_UNCONNECTED_307 VDD VSS DFF_X1 
Xc0_r2_reg_6_ n496 n9_G2B1I1 c0_r2[6] SYNOPSYS_UNCONNECTED_306 VDD VSS DFF_X1 
Xc0_r1_reg_6_ c0[6] n7_G2B1I2 c0_r1[6] SYNOPSYS_UNCONNECTED_305 VDD VSS DFF_X1 
Xc0_r4_reg_7_ n492 n8_G2B1I6 c0_r4[7] SYNOPSYS_UNCONNECTED_304 VDD VSS DFF_X1 
Xc0_r3_reg_7_ n488 n8_G2B1I6 c0_r3[7] SYNOPSYS_UNCONNECTED_303 VDD VSS DFF_X1 
Xc0_r2_reg_7_ n484 n8_G2B1I6 c0_r2[7] SYNOPSYS_UNCONNECTED_302 VDD VSS DFF_X1 
Xc0_r1_reg_7_ c0[7] n8_G2B1I6 c0_r1[7] SYNOPSYS_UNCONNECTED_301 VDD VSS DFF_X1 
Xc0_r4_reg_8_ n480 n7_G2B1I4 c0_r4[8] SYNOPSYS_UNCONNECTED_300 VDD VSS DFF_X1 
Xc0_r3_reg_8_ n476 n7_G2B1I4 c0_r3[8] SYNOPSYS_UNCONNECTED_299 VDD VSS DFF_X1 
XU71 data_in[16] rstn N78 VDD VSS AND2_X1 
XU70 rstn data_in[3] N91 VDD VSS AND2_X1 
XU69 data_in[10] rstn N84 VDD VSS AND2_X1 
XU68 data_in[14] rstn N80 VDD VSS AND2_X1 
XU67 data_in[6] rstn N88 VDD VSS AND2_X1 
XU66 n53 n1110 N600 VDD VSS NAND2_X1 
XU65 n44 n1125 n50 VDD VSS AND2_X1 
XU64 n1133 n7310 N611 VDD VSS NAND2_X1 
XU63 n1010 n910 n810 n54 VDD VSS NOR3_X1 
XU62 rstn n710 n6810 n54 n53 VDD VSS AND4_X1 
XU61 n10921 rstn n6810 n44 VDD VSS AND3_X1 
XU60 n7011 n1096 n44 n45 N74 VDD VSS NAND4_X1 
XU59 n1084 n1127 n52 VDD VSS AND2_X1 
XU58 n1084 n7011 n47 VDD VSS AND2_X1 
XU57 n44 n1127 n1096 n51 VDD VSS AND3_X1 
XU56 N1800 n990 VDD VSS INV_X1 
XU55 n55 n990 n29 n56 N196 VDD VSS OAI22_X1 
XU54 N1790 n1000 VDD VSS INV_X1 
XU53 n55 n1000 n30 n56 N195 VDD VSS OAI22_X1 
XU52 N1780 n1011 VDD VSS INV_X1 
XU51 n55 n1011 n31 n56 N194 VDD VSS OAI22_X1 
XU50 N1770 n1020 VDD VSS INV_X1 
XU49 n55 n1020 n32 n56 N193 VDD VSS OAI22_X1 
XU48 N1760 n1030 VDD VSS INV_X1 
XU47 n55 n1030 n33 n56 N192 VDD VSS OAI22_X1 
XU46 N1750 n1040 VDD VSS INV_X1 
XU45 n55 n1040 n34 n56 N191 VDD VSS OAI22_X1 
XU44 N1740 n1050 VDD VSS INV_X1 
XU43 n55 n1050 n35 n56 N190 VDD VSS OAI22_X1 
XU42 N1730 n1060 VDD VSS INV_X1 
XU41 n55 n1060 n36 n56 N189 VDD VSS OAI22_X1 
XU40 N1720 n1070 VDD VSS INV_X1 
XU39 n55 n1070 n37 n56 N188 VDD VSS OAI22_X1 
XU38 N1710 n1080 VDD VSS INV_X1 
XU37 n55 n1080 n38 n56 N187 VDD VSS OAI22_X1 
XU36 N1700 n1090 VDD VSS INV_X1 
XU35 n55 n1090 n39 n56 N186 VDD VSS OAI22_X1 
XU34 N1690 n1100 VDD VSS INV_X1 
XU33 n55 n1100 n40 n56 N185 VDD VSS OAI22_X1 
XU32 N1680 n1111 VDD VSS INV_X1 
XU31 n55 n1111 n41 n56 N184 VDD VSS OAI22_X1 
XU30 N1670 n1120 VDD VSS INV_X1 
XU29 n55 n1120 n42 n56 N183 VDD VSS OAI22_X1 
XU28 n55 n43 n43 n56 N182 VDD VSS OAI22_X1 
XU25 rstn n12 n56 VDD VSS NAND2_X1 
XU24 sign_r[8] rstn n55 VDD VSS NAND2_X1 
XU23 num_lzd[5] rstn N11000 VDD VSS AND2_X1 
XU22 num_lzd[4] rstn N10 VDD VSS AND2_X1 
XU21 num_lzd[2] rstn N8 VDD VSS AND2_X1 
XU20 num_lzd[3] rstn N900 VDD VSS AND2_X1 
XU19 num_lzd[1] rstn N700 VDD VSS AND2_X1 
XU18 num_lzd[0] rstn N610 VDD VSS AND2_X1 
XU17 n52 n1107 N65 VDD VSS NAND2_X1 
XU16 n52 n1115 N64 VDD VSS NAND2_X1 
XU15 n52 n1119 N63 VDD VSS NAND2_X1 
XU14 n51 n1107 N69 VDD VSS NAND2_X1 
XU13 n51 n1115 N68 VDD VSS NAND2_X1 
XU12 n51 n1119 N67 VDD VSS NAND2_X1 
XU11 n47 n45 N7010 VDD VSS NAND2_X1 
XU10 n51 n45 N66 VDD VSS NAND2_X1 
XU9 n52 n45 N620 VDD VSS NAND2_X1 
XU8 n1107 n47 N73 VDD VSS NAND2_X1 
XU6 n1115 n47 N72 VDD VSS NAND2_X1 
XU5 n1119 n47 N71 VDD VSS NAND2_X1 
XU4 N1810 n980 VDD VSS INV_X1 
XU3 n980 n55 N197 VDD VSS NOR2_X1 
Xdata_out_reg_0_ n166 n9_G2B1I1 data_out[0] SYNOPSYS_UNCONNECTED_298 VDD VSS DFF_X1 
Xdata_out_reg_1_ n462 n9_G2B1I2 data_out[1] SYNOPSYS_UNCONNECTED_297 VDD VSS DFF_X1 
Xdata_out_reg_2_ n456 n7_G2B1I1 data_out[2] SYNOPSYS_UNCONNECTED_296 VDD VSS DFF_X1 
Xdata_out_reg_3_ n139 clk_G1B1I5 data_out[3] SYNOPSYS_UNCONNECTED_295 VDD VSS DFF_X1 
Xdata_out_reg_4_ n1304 n8_G2B1I4 data_out[4] SYNOPSYS_UNCONNECTED_294 VDD VSS DFF_X1 
Xdata_out_reg_5_ n165 n61_G2B1I1 data_out[5] SYNOPSYS_UNCONNECTED_293 VDD VSS DFF_X1 
Xdata_out_reg_6_ n164 n61_G2B1I1 data_out[6] SYNOPSYS_UNCONNECTED_292 VDD VSS DFF_X1 
Xdata_out_reg_7_ n138 n61_G2B1I1 data_out[7] SYNOPSYS_UNCONNECTED_291 VDD VSS DFF_X1 
Xdata_out_reg_8_ n1333 n9_G2B1I1 data_out[8] SYNOPSYS_UNCONNECTED_290 VDD VSS DFF_X1 
Xdata_out_reg_9_ n420 n9_G2B1I1 data_out[9] SYNOPSYS_UNCONNECTED_289 VDD VSS DFF_X1 
Xdata_out_reg_10_ n137 n60 data_out[10] SYNOPSYS_UNCONNECTED_288 VDD VSS DFF_X1 
Xdata_out_reg_11_ n408 n60 data_out[11] SYNOPSYS_UNCONNECTED_287 VDD VSS DFF_X1 
Xdata_out_reg_12_ n162 n60_G2B1I1 data_out[12] SYNOPSYS_UNCONNECTED_286 VDD VSS DFF_X1 
Xdata_out_reg_13_ n400 n2 data_out[13] SYNOPSYS_UNCONNECTED_285 VDD VSS DFF_X1 
Xdata_out_reg_14_ n136 n2_G2B1I3 data_out[14] SYNOPSYS_UNCONNECTED_284 VDD VSS DFF_X1 
Xdata_out_reg_15_ n160 n2_G2B1I3 data_out[15] SYNOPSYS_UNCONNECTED_283 VDD VSS DFF_X1 
Xvalid_out_reg n386 n8_G2B1I4 valid_out SYNOPSYS_UNCONNECTED_282 VDD VSS DFF_X1 
Xsum2_rnd_reg_0_ n158 n7 SYNOPSYS_UNCONNECTED_281 n43 VDD VSS DFF_X1 
Xsum2_rnd_reg_1_ n157 n9_G2B1I2 SYNOPSYS_UNCONNECTED_280 n42 VDD VSS DFF_X1 
Xsum2_rnd_reg_2_ n156 n9_G2B1I2 SYNOPSYS_UNCONNECTED_279 n41 VDD VSS DFF_X1 
Xsum2_rnd_reg_3_ n155 n9_G2B1I2 SYNOPSYS_UNCONNECTED_278 n40 VDD VSS DFF_X1 
Xsum2_rnd_reg_4_ n154 n7_G2B1I2 SYNOPSYS_UNCONNECTED_277 n39 VDD VSS DFF_X1 
Xsum2_rnd_reg_5_ n153 n7 SYNOPSYS_UNCONNECTED_276 n38 VDD VSS DFF_X1 
Xsum2_rnd_reg_6_ n152 n7 SYNOPSYS_UNCONNECTED_275 n37 VDD VSS DFF_X1 
Xsum2_rnd_reg_7_ n151 n62 SYNOPSYS_UNCONNECTED_274 n36 VDD VSS DFF_X1 
XU141 sum2[8] n5 n940 VDD VSS XOR2_X1 
XU140 sum2[7] n17 n930 VDD VSS XOR2_X1 
XU139 sum2[6] n16 n920 VDD VSS XOR2_X1 
XU138 sum2[5] n4 n911 VDD VSS XOR2_X1 
XU137 sum2[4] n3 n9000 VDD VSS XOR2_X1 
XU136 sum2[2] sum2[3] n890 VDD VSS XOR2_X1 
XU135 n870 n880 N92 VDD VSS NOR2_X1 
XU134 n850 n860 N93 VDD VSS NOR2_X1 
XU133 n830 n840 N94 VDD VSS NOR2_X1 
XU132 n811 n820 N95 VDD VSS NOR2_X1 
XU131 n790 n800 N96 VDD VSS NOR2_X1 
XU130 n770 n780 N97 VDD VSS NOR2_X1 
XU129 n750 n760 N98 VDD VSS NOR2_X1 
XU128 n730 n740 N99 VDD VSS NOR2_X1 
XU127 n711 n720 N100 VDD VSS NOR2_X1 
XU126 n690 n7000 N101 VDD VSS NOR2_X1 
XU125 n670 n680 N102 VDD VSS NOR2_X1 
XU124 n650 n660 N103 VDD VSS NOR2_X1 
XU123 n630 n640 N104 VDD VSS NOR2_X1 
XU122 n6110 n6200 N105 VDD VSS NOR2_X1 
XU121 n59 n6000 N106 VDD VSS NOR2_X1 
XU120 n1091 n1095 n46 VDD VSS NOR2_X1 
XU119 n1091 n7310 n48 VDD VSS NOR2_X1 
XU118 n1095 n7210 n49 VDD VSS NOR2_X1 
XU117 n1086 n7310 n45 VDD VSS NOR2_X1 
XU116 sum2[16] n15 n950 VDD VSS NAND2_X1 
XU115 n58 n950 n57 VDD VSS XOR2_X1 
XU114 sum2[16] n15 n28 VDD VSS XOR2_X1 
XU113 sum2[15] n21 n27 VDD VSS XOR2_X1 
XU112 sum2[14] n20 n26 VDD VSS XOR2_X1 
XU111 sum2[13] n14 n25 VDD VSS XOR2_X1 
XU110 sum2[12] n19 n24 VDD VSS XOR2_X1 
XU109 sum2[11] n18 n23 VDD VSS XOR2_X1 
XU108 sum2[10] n13 n22 VDD VSS XOR2_X1 
XU107 sum2[14] n20 n21 VDD VSS AND2_X1 
XU106 sum2[13] n14 n20 VDD VSS AND2_X1 
XU105 sum2[11] n18 n19 VDD VSS AND2_X1 
XU104 sum2[10] n13 n18 VDD VSS AND2_X1 
XU103 sum2[6] n16 n17 VDD VSS AND2_X1 
XU102 sum2[5] n4 n16 VDD VSS AND2_X1 
XU101 sum2[15] n21 n15 VDD VSS AND2_X1 
XU100 sum2[12] n19 n14 VDD VSS AND2_X1 
XU99 sum2[9] n6100 n13 VDD VSS AND2_X1 
XU98 sum2[8] n5 n6100 VDD VSS AND2_X1 
XU97 sum2[7] n17 n5 VDD VSS AND2_X1 
XU96 sum2[4] n3 n4 VDD VSS AND2_X1 
XU95 sum2[2] sum2[3] n3 VDD VSS AND2_X1 
XU94 sum2[9] n6100 n1 VDD VSS XOR2_X1 
XU93 data_in[1] IN1 N76 VDD VSS AND2_X1 
XU92 data_in[2] IN0 N75 VDD VSS AND2_X1 
XU91 data_in[17] rstn N77 VDD VSS AND2_X1 
XU90 valid_in IN2 N107 VDD VSS AND2_X1 
XU89 valid_in_r[0] IN2 N108 VDD VSS AND2_X1 
XU88 n704 IN1 N109 VDD VSS AND2_X1 
XU87 valid_in_r[2] IN1 N11010 VDD VSS AND2_X1 
XU86 valid_in_r[3] IN1 N111 VDD VSS AND2_X1 
XU85 valid_in_r[4] IN1 N112 VDD VSS AND2_X1 
XU84 valid_in_r[5] IN1 N113 VDD VSS AND2_X1 
XU83 valid_in_r[6] IN1 N114 VDD VSS AND2_X1 
XU82 valid_in_r[7] IN1 N115 VDD VSS AND2_X1 
XU81 valid_in_r[8] IN1 N147 VDD VSS AND2_X1 
XU80 data_in[4] rstn N9010 VDD VSS AND2_X1 
XU79 data_in[5] rstn N89 VDD VSS AND2_X1 
XU78 data_in[7] rstn N87 VDD VSS AND2_X1 
XU77 data_in[8] rstn N86 VDD VSS AND2_X1 
XU76 data_in[9] rstn N85 VDD VSS AND2_X1 
XU75 data_in[11] rstn N83 VDD VSS AND2_X1 
XU74 data_in[12] rstn N82 VDD VSS AND2_X1 
XU73 data_in[13] rstn N81 VDD VSS AND2_X1 
XU72 data_in[15] rstn N79 VDD VSS AND2_X1 
XU145 clk_G1B1I7 n6111 VDD VSS BUF_X32 
XU142 clk_G1B1I7 n10920 VDD VSS BUF_X32 
XCLKBUF_X1_G2B1I1 n11 n11_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I2 n11 n11_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I3 n11 n11_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I4 n11 n11_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I5 n11 n11_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I6 n11 n11_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I7 n11 n11_G2B1I7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I31 n2 n2_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I13 n10920 n10_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I23 n10920 n10_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I33 n10920 n10_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I42 n10920 n10_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I25 n6310 n63_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I15 clk_G1B1I5 n8_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I26 clk_G1B1I5 n8_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I44 clk_G1B1I5 n8_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I53 clk_G1B1I5 n8_G2B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I61 clk_G1B1I5 n8_G2B1I6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I71 clk_G1B1I5 n8_G2B1I7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I81 clk_G1B1I5 n8_G2B1I8 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I16 n7 n7_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I27 n7 n7_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I45 n7 n7_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I29 n62 n62_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I19 n6111 n61_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X3_G1B1I7 clk clk_G1B1I7 VDD VSS CLKBUF_X3 
XCLKBUF_X3_G1B1I8 clk clk_G1B1I8 VDD VSS CLKBUF_X1 
XCLKBUF_X2_G1B1I5 clk clk_G1B1I5 VDD VSS CLKBUF_X1 
XCLKBUF_X3_G1B1I4 clk clk_G1B1I4 VDD VSS CLKBUF_X1 
XU146 clk_G1B1I4 n62 VDD VSS CLKBUF_X1 
XU27 clk_G1B1I4 n9 VDD VSS CLKBUF_X1 
XCLKBUF_X2_G1B1I1 clk clk_G1B1I1 VDD VSS CLKBUF_X1 
XU1 clk_cts_3 n2 VDD VSS CLKBUF_X1 
XU143 clk_cts_3 n11 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I8 n6310 n63_G2B1I8 VDD VSS CLKBUF_X1 
XU7 clk_G1B1I4 n7 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I17 n9 n9_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I28 n9 n9_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I22 n6 n6_G2B1I2 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I32 n6 n6_G2B1I3 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I41 n6 n6_G2B1I4 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I51 n6 n6_G2B1I5 VDD VSS CLKBUF_X1 
XU2 clk_G1B1I8 n6 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I14 n60 n60_G2B1I1 VDD VSS CLKBUF_X1 
XCLKBUF_X1_G2B1I52 n60 n60_G2B1I5 VDD VSS CLKBUF_X1 
XU144 clk_G1B1I8 n60 VDD VSS CLKBUF_X1 
XU147 clk_G1B1I1 n6310 VDD VSS CLKBUF_X3 
XU26 num_lzd_r[0] n132 VDD VSS CLKBUF_X2 
XU149 n204 n133 VDD VSS BUF_X1 
XU151 n1101 n134 VDD VSS BUF_X1 
XU154 n208 n135 VDD VSS BUF_X1 
XU155 n161 n136 VDD VSS BUF_X1 
XU156 n415 n137 VDD VSS BUF_X1 
XU157 n163 n138 VDD VSS BUF_X1 
XU158 n452 n139 VDD VSS BUF_X1 
XU159 n589 n140 VDD VSS BUF_X1 
XU160 n866 n141 VDD VSS BUF_X1 
XU161 n1088 n142 VDD VSS BUF_X1 
XU162 num_lzd_r[2] n143 VDD VSS BUF_X1 
XU163 n1123 n1127 VDD VSS INV_X16 
XU164 n1116 n1117 VDD VSS INV_X8 
XU165 n1108 n1109 VDD VSS INV_X1 
XU166 n1102 n1103 VDD VSS INV_X1 
XU167 n1890 n1900 VDD VSS INV_X1 
XU168 n144 n145 VDD VSS INV_X4 
XU169 n146 n1470 VDD VSS INV_X4 
XU170 n149 n150 VDD VSS INV_X1 
XU171 n238 n144 VDD VSS INV_X1 
XU172 n254 n146 VDD VSS INV_X1 
XU173 n274 n148 VDD VSS BUF_X1 
XU174 n273 n149 VDD VSS INV_X1 
XU175 n347 n151 VDD VSS BUF_X1 
XU176 n350 n152 VDD VSS BUF_X1 
XU177 n357 n153 VDD VSS BUF_X1 
XU178 n362 n154 VDD VSS BUF_X1 
XU179 n367 n155 VDD VSS BUF_X1 
XU180 n372 n156 VDD VSS BUF_X1 
XU181 n377 n157 VDD VSS BUF_X1 
XU182 n382 n158 VDD VSS BUF_X1 
XU183 n389 n159 VDD VSS INV_X1 
XU184 n159 n160 VDD VSS INV_X8 
XU185 n395 n161 VDD VSS CLKBUF_X1 
XU186 n407 n162 VDD VSS BUF_X1 
XU187 n431 n163 VDD VSS CLKBUF_X1 
XU188 n437 n164 VDD VSS BUF_X1 
XU189 n443 n165 VDD VSS BUF_X1 
XU190 n470 n166 VDD VSS BUF_X1 
XU191 n737 n167 VDD VSS BUF_X1 
XU192 n743 n168 VDD VSS BUF_X1 
XU193 n748 n169 VDD VSS BUF_X1 
XU194 n754 n170 VDD VSS BUF_X1 
XU195 n765 n171 VDD VSS CLKBUF_X1 
XU196 n771 n172 VDD VSS INV_X1 
XU197 n172 n173 VDD VSS INV_X8 
XU198 n778 n174 VDD VSS INV_X1 
XU199 n174 n175 VDD VSS INV_X16 
XU200 n795 n176 VDD VSS BUF_X1 
XU201 n809 n177 VDD VSS INV_X1 
XU202 n177 n178 VDD VSS INV_X16 
XU203 n825 n179 VDD VSS INV_X1 
XU204 n179 n180 VDD VSS INV_X16 
XU205 n834 n181 VDD VSS BUF_X1 
XU206 n838 n1820 VDD VSS BUF_X1 
XU207 n855 n1830 VDD VSS INV_X1 
XU208 n1830 n1840 VDD VSS INV_X16 
XU209 n921 n1850 VDD VSS BUF_X1 
XU210 n929 n1860 VDD VSS BUF_X1 
XU211 n1017 n1870 VDD VSS CLKBUF_X1 
XU212 n1057 n1880 VDD VSS BUF_X1 
XU213 n1056 n1890 VDD VSS INV_X1 
XU214 N610 n1910 VDD VSS INV_X1 
XU215 n1910 n1920 VDD VSS INV_X16 
XU216 n1158 n1930 VDD VSS CLKBUF_X1 
XU217 n1202 n1940 VDD VSS BUF_X1 
XU218 n1216 n1950 VDD VSS BUF_X1 
XU219 n1229 n1960 VDD VSS INV_X1 
XU220 n1960 n1970 VDD VSS INV_X16 
XU221 n1245 n198 VDD VSS BUF_X1 
XU222 n1258 n199 VDD VSS INV_X1 
XU223 n199 n200 VDD VSS INV_X16 
XU224 n1299 n201 VDD VSS BUF_X1 
XU225 offset[1] n202 VDD VSS CLKBUF_X1 
XU226 num_lzd_r[1] n203 VDD VSS INV_X1 
XU227 n203 n204 VDD VSS INV_X32 
XU228 n134 n205 VDD VSS BUF_X1 
XU229 offset[0] n206 VDD VSS INV_X32 
XU230 n206 n207 VDD VSS INV_X1 
XU231 n1098 n208 VDD VSS BUF_X1 
XU232 n1289 n209 VDD VSS BUF_X1 
XU233 n799 n210 VDD VSS BUF_X1 
XU234 c1_r1[17] n211 VDD VSS CLKBUF_X1 
XU235 n213 n212 VDD VSS CLKBUF_X1 
XU236 n211 n213 VDD VSS INV_X32 
XU237 n212 n214 VDD VSS INV_X32 
XU238 c1_r1[16] n215 VDD VSS CLKBUF_X1 
XU239 n217 n216 VDD VSS CLKBUF_X1 
XU240 n215 n217 VDD VSS INV_X32 
XU241 n216 n218 VDD VSS INV_X32 
XU242 c1_r1[15] n219 VDD VSS CLKBUF_X1 
XU243 n221 n220 VDD VSS CLKBUF_X1 
XU244 n219 n221 VDD VSS INV_X32 
XU245 n220 n222 VDD VSS INV_X32 
XU246 c1_r1[14] n223 VDD VSS CLKBUF_X1 
XU247 n225 n224 VDD VSS CLKBUF_X1 
XU248 n223 n225 VDD VSS INV_X32 
XU249 n224 n226 VDD VSS INV_X32 
XU250 c1_r1[13] n227 VDD VSS CLKBUF_X1 
XU251 n229 n228 VDD VSS CLKBUF_X1 
XU252 n227 n229 VDD VSS INV_X32 
XU253 n228 n230 VDD VSS INV_X32 
XU254 c1_r1[12] n231 VDD VSS CLKBUF_X1 
XU255 n233 n232 VDD VSS CLKBUF_X1 
XU256 n231 n233 VDD VSS INV_X32 
XU257 n232 n234 VDD VSS INV_X32 
XU258 c1_r1[11] n235 VDD VSS CLKBUF_X1 
XU259 n237 n236 VDD VSS CLKBUF_X1 
XU260 n235 n237 VDD VSS INV_X32 
XU261 n236 n238 VDD VSS INV_X32 
XU262 c1_r1[10] n239 VDD VSS CLKBUF_X1 
XU263 n241 n240 VDD VSS CLKBUF_X1 
XU264 n239 n241 VDD VSS INV_X32 
XU265 n240 n242 VDD VSS INV_X32 
XU266 c1_r1[9] n243 VDD VSS CLKBUF_X1 
XU267 n245 n244 VDD VSS CLKBUF_X1 
XU268 n243 n245 VDD VSS INV_X32 
XU269 n244 n246 VDD VSS INV_X32 
XU270 c1_r1[8] n247 VDD VSS CLKBUF_X1 
XU271 n249 n248 VDD VSS CLKBUF_X1 
XU272 n247 n249 VDD VSS INV_X32 
XU273 n248 n250 VDD VSS INV_X32 
XU274 c1_r1[7] n251 VDD VSS CLKBUF_X1 
XU275 n253 n252 VDD VSS CLKBUF_X1 
XU276 n251 n253 VDD VSS INV_X32 
XU277 n252 n254 VDD VSS INV_X32 
XU278 c1_r1[6] n255 VDD VSS CLKBUF_X1 
XU279 n257 n256 VDD VSS CLKBUF_X1 
XU280 n255 n257 VDD VSS INV_X32 
XU281 n256 n258 VDD VSS INV_X32 
XU282 c1_r1[5] n259 VDD VSS CLKBUF_X1 
XU283 n261 n260 VDD VSS CLKBUF_X1 
XU284 n259 n261 VDD VSS INV_X32 
XU285 n260 n262 VDD VSS INV_X32 
XU286 c1_r1[4] n263 VDD VSS CLKBUF_X1 
XU287 n265 n264 VDD VSS CLKBUF_X1 
XU288 n263 n265 VDD VSS INV_X32 
XU289 n264 n266 VDD VSS INV_X32 
XU290 c1_r1[3] n267 VDD VSS CLKBUF_X1 
XU291 n269 n268 VDD VSS CLKBUF_X1 
XU292 n267 n269 VDD VSS INV_X32 
XU293 n268 n270 VDD VSS INV_X32 
XU294 c1_r1[2] n271 VDD VSS CLKBUF_X1 
XU295 n150 n272 VDD VSS CLKBUF_X1 
XU296 n271 n273 VDD VSS INV_X32 
XU297 n272 n274 VDD VSS INV_X32 
XU298 c1_r1[1] n275 VDD VSS CLKBUF_X1 
XU299 n277 n276 VDD VSS CLKBUF_X1 
XU300 n275 n277 VDD VSS INV_X32 
XU301 n276 n278 VDD VSS INV_X32 
XU302 c1_r1[0] n279 VDD VSS CLKBUF_X1 
XU303 n281 n280 VDD VSS CLKBUF_X1 
XU304 n279 n281 VDD VSS INV_X32 
XU305 n280 n282 VDD VSS INV_X32 
XU306 x_r4[14] n283 VDD VSS CLKBUF_X1 
XU307 n285 n284 VDD VSS CLKBUF_X1 
XU308 n283 n285 VDD VSS INV_X32 
XU309 n284 n286 VDD VSS INV_X32 
XU310 x_r4[13] n287 VDD VSS CLKBUF_X1 
XU311 n289 n288 VDD VSS CLKBUF_X1 
XU312 n287 n289 VDD VSS INV_X32 
XU313 n288 n290 VDD VSS INV_X32 
XU314 x_r4[12] n291 VDD VSS CLKBUF_X1 
XU315 n293 n292 VDD VSS CLKBUF_X1 
XU316 n291 n293 VDD VSS INV_X32 
XU317 n292 n294 VDD VSS INV_X32 
XU318 x_r4[11] n295 VDD VSS CLKBUF_X1 
XU319 n297 n296 VDD VSS CLKBUF_X1 
XU320 n295 n297 VDD VSS INV_X32 
XU321 n296 n298 VDD VSS INV_X32 
XU322 x_r4[10] n299 VDD VSS CLKBUF_X1 
XU323 n301 n300 VDD VSS CLKBUF_X1 
XU324 n299 n301 VDD VSS INV_X32 
XU325 n300 n302 VDD VSS INV_X32 
XU326 x_r4[9] n303 VDD VSS CLKBUF_X1 
XU327 n305 n304 VDD VSS CLKBUF_X1 
XU328 n303 n305 VDD VSS INV_X32 
XU329 n304 n306 VDD VSS INV_X32 
XU330 x_r4[8] n307 VDD VSS CLKBUF_X1 
XU331 n309 n308 VDD VSS CLKBUF_X1 
XU332 n307 n309 VDD VSS INV_X32 
XU333 n308 n310 VDD VSS INV_X32 
XU334 x_r4[7] n311 VDD VSS CLKBUF_X1 
XU335 n313 n312 VDD VSS CLKBUF_X1 
XU336 n311 n313 VDD VSS INV_X32 
XU337 n312 n314 VDD VSS INV_X32 
XU338 x_r4[6] n315 VDD VSS CLKBUF_X1 
XU339 n317 n316 VDD VSS CLKBUF_X1 
XU340 n315 n317 VDD VSS INV_X32 
XU341 n316 n318 VDD VSS INV_X32 
XU342 x_r4[5] n319 VDD VSS CLKBUF_X1 
XU343 n321 n320 VDD VSS CLKBUF_X1 
XU344 n319 n321 VDD VSS INV_X32 
XU345 n320 n322 VDD VSS INV_X32 
XU346 x_r4[4] n323 VDD VSS CLKBUF_X1 
XU347 n325 n324 VDD VSS CLKBUF_X1 
XU348 n323 n325 VDD VSS INV_X32 
XU349 n324 n326 VDD VSS INV_X32 
XU350 x_r4[3] n327 VDD VSS CLKBUF_X1 
XU351 n329 n328 VDD VSS CLKBUF_X1 
XU352 n327 n329 VDD VSS INV_X32 
XU353 n328 n330 VDD VSS INV_X32 
XU354 x_r4[2] n331 VDD VSS CLKBUF_X1 
XU355 n333 n332 VDD VSS CLKBUF_X1 
XU356 n331 n333 VDD VSS INV_X32 
XU357 n332 n334 VDD VSS INV_X32 
XU358 x_r4[1] n335 VDD VSS CLKBUF_X1 
XU359 n337 n336 VDD VSS CLKBUF_X1 
XU360 n335 n337 VDD VSS INV_X32 
XU361 n336 n338 VDD VSS INV_X32 
XU362 x_r4[0] n339 VDD VSS CLKBUF_X1 
XU363 n341 n340 VDD VSS CLKBUF_X1 
XU364 n339 n341 VDD VSS INV_X32 
XU365 n340 n342 VDD VSS INV_X32 
XU366 n346 n343 VDD VSS CLKBUF_X1 
XU367 n343 n344 VDD VSS INV_X32 
XU368 n344 n345 VDD VSS INV_X1 
XU369 n22 n346 VDD VSS INV_X1 
XU370 n345 n347 VDD VSS INV_X32 
XU371 n349 n348 VDD VSS CLKBUF_X1 
XU372 n352 n349 VDD VSS INV_X1 
XU373 n348 n350 VDD VSS INV_X32 
XU374 n1 n351 VDD VSS INV_X1 
XU375 n351 n352 VDD VSS INV_X32 
XU376 n356 n353 VDD VSS CLKBUF_X1 
XU377 n353 n354 VDD VSS INV_X32 
XU378 n354 n355 VDD VSS INV_X1 
XU379 n940 n356 VDD VSS INV_X1 
XU380 n355 n357 VDD VSS INV_X32 
XU381 n361 n358 VDD VSS CLKBUF_X1 
XU382 n358 n359 VDD VSS INV_X32 
XU383 n359 n360 VDD VSS INV_X1 
XU384 n930 n361 VDD VSS INV_X1 
XU385 n360 n362 VDD VSS INV_X32 
XU386 n366 n363 VDD VSS CLKBUF_X1 
XU387 n363 n364 VDD VSS INV_X32 
XU388 n364 n365 VDD VSS INV_X1 
XU389 n920 n366 VDD VSS INV_X1 
XU390 n365 n367 VDD VSS INV_X32 
XU391 n371 n368 VDD VSS CLKBUF_X1 
XU392 n368 n369 VDD VSS INV_X32 
XU393 n369 n370 VDD VSS INV_X1 
XU394 n911 n371 VDD VSS INV_X1 
XU395 n370 n372 VDD VSS INV_X32 
XU396 n376 n373 VDD VSS CLKBUF_X1 
XU397 n373 n374 VDD VSS INV_X32 
XU398 n374 n375 VDD VSS INV_X1 
XU399 n9000 n376 VDD VSS INV_X1 
XU400 n375 n377 VDD VSS INV_X32 
XU401 n381 n378 VDD VSS CLKBUF_X1 
XU402 n378 n379 VDD VSS INV_X32 
XU403 n379 n380 VDD VSS INV_X1 
XU404 n890 n381 VDD VSS INV_X1 
XU405 n380 n382 VDD VSS INV_X32 
XU406 N147 n383 VDD VSS CLKBUF_X1 
XU407 n385 n384 VDD VSS CLKBUF_X1 
XU408 n383 n385 VDD VSS INV_X32 
XU409 n384 n386 VDD VSS INV_X32 
XU410 n388 n387 VDD VSS CLKBUF_X1 
XU411 n391 n388 VDD VSS INV_X1 
XU412 n387 n389 VDD VSS INV_X32 
XU413 N197 n390 VDD VSS INV_X1 
XU414 n390 n391 VDD VSS INV_X32 
XU415 n394 n392 VDD VSS INV_X32 
XU416 n392 n393 VDD VSS INV_X1 
XU417 n397 n394 VDD VSS INV_X1 
XU418 n393 n395 VDD VSS INV_X32 
XU419 N196 n396 VDD VSS INV_X1 
XU420 n396 n397 VDD VSS INV_X32 
XU421 n399 n398 VDD VSS CLKBUF_X1 
XU422 n402 n399 VDD VSS INV_X1 
XU423 n398 n400 VDD VSS INV_X32 
XU424 N195 n401 VDD VSS INV_X1 
XU425 n401 n402 VDD VSS INV_X32 
XU426 n405 n403 VDD VSS CLKBUF_X1 
XU427 n406 n404 VDD VSS INV_X32 
XU428 n404 n405 VDD VSS INV_X1 
XU429 N194 n406 VDD VSS INV_X1 
XU430 n403 n407 VDD VSS INV_X32 
XU431 n410 n408 VDD VSS CLKBUF_X1 
XU432 n412 n409 VDD VSS INV_X1 
XU433 n409 n410 VDD VSS INV_X32 
XU434 N193 n411 VDD VSS INV_X1 
XU435 n411 n412 VDD VSS INV_X32 
XU436 N192 n413 VDD VSS BUF_X16 
XU437 n417 n414 VDD VSS INV_X1 
XU438 n414 n415 VDD VSS INV_X32 
XU439 n413 n416 VDD VSS INV_X1 
XU440 n416 n417 VDD VSS INV_X32 
XU441 n419 n418 VDD VSS CLKBUF_X1 
XU442 n422 n419 VDD VSS INV_X1 
XU443 n418 n420 VDD VSS INV_X32 
XU444 N191 n421 VDD VSS INV_X1 
XU445 n421 n422 VDD VSS INV_X32 
XU446 n424 n423 VDD VSS CLKBUF_X1 
XU447 n427 n424 VDD VSS INV_X1 
XU448 n423 n425 VDD VSS INV_X32 
XU449 N190 n426 VDD VSS INV_X1 
XU450 n426 n427 VDD VSS INV_X32 
XU451 n430 n428 VDD VSS INV_X32 
XU452 n428 n429 VDD VSS INV_X1 
XU453 n433 n430 VDD VSS INV_X1 
XU454 n429 n431 VDD VSS INV_X32 
XU455 N189 n432 VDD VSS INV_X1 
XU456 n432 n433 VDD VSS INV_X32 
XU457 n436 n434 VDD VSS INV_X32 
XU458 n434 n435 VDD VSS INV_X1 
XU459 n439 n436 VDD VSS INV_X1 
XU460 n435 n437 VDD VSS INV_X32 
XU461 N188 n438 VDD VSS INV_X1 
XU462 n438 n439 VDD VSS INV_X32 
XU463 n442 n440 VDD VSS INV_X32 
XU464 n440 n441 VDD VSS INV_X1 
XU465 n445 n442 VDD VSS INV_X1 
XU466 n441 n443 VDD VSS INV_X32 
XU467 N187 n444 VDD VSS INV_X1 
XU468 n444 n445 VDD VSS INV_X32 
XU469 n448 n446 VDD VSS CLKBUF_X1 
XU470 n450 n447 VDD VSS INV_X1 
XU471 n447 n448 VDD VSS INV_X32 
XU472 N186 n449 VDD VSS INV_X1 
XU473 n449 n450 VDD VSS INV_X32 
XU474 n454 n451 VDD VSS INV_X1 
XU475 n451 n452 VDD VSS INV_X32 
XU476 N185 n453 VDD VSS INV_X1 
XU477 n453 n454 VDD VSS INV_X32 
XU478 n458 n455 VDD VSS INV_X1 
XU479 n455 n456 VDD VSS INV_X32 
XU480 n460 n457 VDD VSS INV_X1 
XU481 n457 n458 VDD VSS INV_X32 
XU482 N184 n459 VDD VSS INV_X1 
XU483 n459 n460 VDD VSS INV_X32 
XU484 n464 n461 VDD VSS INV_X1 
XU485 n461 n462 VDD VSS INV_X32 
XU486 n466 n463 VDD VSS INV_X1 
XU487 n463 n464 VDD VSS INV_X32 
XU488 N183 n465 VDD VSS INV_X1 
XU489 n465 n466 VDD VSS INV_X32 
XU490 n469 n467 VDD VSS INV_X32 
XU491 n467 n468 VDD VSS INV_X1 
XU492 n472 n469 VDD VSS INV_X1 
XU493 n468 n470 VDD VSS INV_X32 
XU494 N182 n471 VDD VSS INV_X1 
XU495 n471 n472 VDD VSS INV_X32 
XU496 c0_r2[8] n473 VDD VSS CLKBUF_X1 
XU497 n475 n474 VDD VSS CLKBUF_X1 
XU498 n473 n475 VDD VSS INV_X32 
XU499 n474 n476 VDD VSS INV_X32 
XU500 c0_r3[8] n477 VDD VSS CLKBUF_X1 
XU501 n479 n478 VDD VSS CLKBUF_X1 
XU502 n477 n479 VDD VSS INV_X32 
XU503 n478 n480 VDD VSS INV_X32 
XU504 c0_r1[7] n481 VDD VSS CLKBUF_X1 
XU505 n483 n482 VDD VSS CLKBUF_X1 
XU506 n481 n483 VDD VSS INV_X32 
XU507 n482 n484 VDD VSS INV_X32 
XU508 c0_r2[7] n485 VDD VSS CLKBUF_X1 
XU509 n487 n486 VDD VSS CLKBUF_X1 
XU510 n485 n487 VDD VSS INV_X32 
XU511 n486 n488 VDD VSS INV_X32 
XU512 c0_r3[7] n489 VDD VSS CLKBUF_X1 
XU513 n491 n490 VDD VSS CLKBUF_X1 
XU514 n489 n491 VDD VSS INV_X32 
XU515 n490 n492 VDD VSS INV_X32 
XU516 c0_r1[6] n493 VDD VSS CLKBUF_X1 
XU517 n495 n494 VDD VSS CLKBUF_X1 
XU518 n493 n495 VDD VSS INV_X32 
XU519 n494 n496 VDD VSS INV_X32 
XU520 c0_r2[6] n497 VDD VSS CLKBUF_X1 
XU521 n499 n498 VDD VSS CLKBUF_X1 
XU522 n497 n499 VDD VSS INV_X32 
XU523 n498 n500 VDD VSS INV_X32 
XU524 c0_r3[6] n501 VDD VSS CLKBUF_X1 
XU525 n503 n502 VDD VSS CLKBUF_X1 
XU526 n501 n503 VDD VSS INV_X32 
XU527 n502 n504 VDD VSS INV_X32 
XU528 c0_r1[5] n505 VDD VSS CLKBUF_X1 
XU529 n507 n506 VDD VSS CLKBUF_X1 
XU530 n505 n507 VDD VSS INV_X32 
XU531 n506 n508 VDD VSS INV_X32 
XU532 c0_r2[5] n509 VDD VSS CLKBUF_X1 
XU533 n511 n510 VDD VSS CLKBUF_X1 
XU534 n509 n511 VDD VSS INV_X32 
XU535 n510 n512 VDD VSS INV_X32 
XU536 c0_r3[5] n513 VDD VSS CLKBUF_X1 
XU537 n515 n514 VDD VSS CLKBUF_X1 
XU538 n513 n515 VDD VSS INV_X32 
XU539 n514 n516 VDD VSS INV_X32 
XU540 c0_r1[4] n517 VDD VSS CLKBUF_X1 
XU541 n519 n518 VDD VSS CLKBUF_X1 
XU542 n517 n519 VDD VSS INV_X32 
XU543 n518 n520 VDD VSS INV_X32 
XU544 c0_r2[4] n521 VDD VSS CLKBUF_X1 
XU545 n523 n522 VDD VSS CLKBUF_X1 
XU546 n521 n523 VDD VSS INV_X32 
XU547 n522 n524 VDD VSS INV_X32 
XU548 c0_r3[4] n525 VDD VSS CLKBUF_X1 
XU549 n527 n526 VDD VSS CLKBUF_X1 
XU550 n525 n527 VDD VSS INV_X32 
XU551 n526 n528 VDD VSS INV_X32 
XU552 c0_r1[3] n529 VDD VSS CLKBUF_X1 
XU553 n531 n530 VDD VSS CLKBUF_X1 
XU554 n529 n531 VDD VSS INV_X32 
XU555 n530 n532 VDD VSS INV_X32 
XU556 c0_r2[3] n533 VDD VSS CLKBUF_X1 
XU557 n535 n534 VDD VSS CLKBUF_X1 
XU558 n533 n535 VDD VSS INV_X32 
XU559 n534 n536 VDD VSS INV_X32 
XU560 c0_r3[3] n537 VDD VSS CLKBUF_X1 
XU561 n539 n538 VDD VSS CLKBUF_X1 
XU562 n537 n539 VDD VSS INV_X32 
XU563 n538 n540 VDD VSS INV_X32 
XU564 c0_r1[2] n541 VDD VSS CLKBUF_X1 
XU565 n543 n542 VDD VSS CLKBUF_X1 
XU566 n541 n543 VDD VSS INV_X32 
XU567 n542 n544 VDD VSS INV_X32 
XU568 c0_r2[2] n545 VDD VSS CLKBUF_X1 
XU569 n547 n546 VDD VSS CLKBUF_X1 
XU570 n545 n547 VDD VSS INV_X32 
XU571 n546 n548 VDD VSS INV_X32 
XU572 c0_r3[2] n549 VDD VSS CLKBUF_X1 
XU573 n551 n550 VDD VSS CLKBUF_X1 
XU574 n549 n551 VDD VSS INV_X32 
XU575 n550 n552 VDD VSS INV_X32 
XU576 c0_r1[1] n553 VDD VSS CLKBUF_X1 
XU577 n555 n554 VDD VSS CLKBUF_X1 
XU578 n553 n555 VDD VSS INV_X32 
XU579 n554 n556 VDD VSS INV_X32 
XU580 c0_r2[1] n557 VDD VSS CLKBUF_X1 
XU581 n559 n558 VDD VSS CLKBUF_X1 
XU582 n557 n559 VDD VSS INV_X32 
XU583 n558 n560 VDD VSS INV_X32 
XU584 c0_r3[1] n561 VDD VSS CLKBUF_X1 
XU585 n563 n562 VDD VSS CLKBUF_X1 
XU586 n561 n563 VDD VSS INV_X32 
XU587 n562 n564 VDD VSS INV_X32 
XU588 c0_r1[0] n565 VDD VSS CLKBUF_X1 
XU589 n567 n566 VDD VSS CLKBUF_X1 
XU590 n565 n567 VDD VSS INV_X32 
XU591 n566 n568 VDD VSS INV_X32 
XU592 c0_r2[0] n569 VDD VSS CLKBUF_X1 
XU593 n571 n570 VDD VSS CLKBUF_X1 
XU594 n569 n571 VDD VSS INV_X32 
XU595 n570 n572 VDD VSS INV_X32 
XU596 c0_r3[0] n573 VDD VSS CLKBUF_X1 
XU597 n575 n574 VDD VSS CLKBUF_X1 
XU598 n573 n575 VDD VSS INV_X32 
XU599 n574 n576 VDD VSS INV_X32 
XU600 c0_r4[17] n577 VDD VSS CLKBUF_X1 
XU601 n579 n578 VDD VSS CLKBUF_X1 
XU602 n577 n579 VDD VSS INV_X32 
XU603 n578 n580 VDD VSS INV_X32 
XU604 c0_r4[16] n581 VDD VSS CLKBUF_X1 
XU605 n583 n582 VDD VSS CLKBUF_X1 
XU606 n581 n583 VDD VSS INV_X32 
XU607 n582 n584 VDD VSS INV_X32 
XU608 c0_r4[15] n585 VDD VSS CLKBUF_X1 
XU609 n587 n586 VDD VSS CLKBUF_X1 
XU610 n585 n587 VDD VSS INV_X32 
XU611 n586 n588 VDD VSS INV_X32 
XU612 n592 n589 VDD VSS CLKBUF_X1 
XU613 n591 n590 VDD VSS CLKBUF_X1 
XU614 c0_r4[14] n591 VDD VSS INV_X32 
XU615 n590 n592 VDD VSS INV_X32 
XU616 c0_r4[13] n593 VDD VSS CLKBUF_X1 
XU617 n595 n594 VDD VSS CLKBUF_X1 
XU618 n593 n595 VDD VSS INV_X32 
XU619 n594 n596 VDD VSS INV_X32 
XU620 c0_r4[12] n597 VDD VSS CLKBUF_X1 
XU621 n599 n598 VDD VSS CLKBUF_X1 
XU622 n597 n599 VDD VSS INV_X32 
XU623 n598 n601 VDD VSS INV_X32 
XU624 c0_r4[11] n602 VDD VSS CLKBUF_X1 
XU625 n604 n603 VDD VSS CLKBUF_X1 
XU626 n602 n604 VDD VSS INV_X32 
XU627 n603 n605 VDD VSS INV_X32 
XU628 c0_r4[10] n606 VDD VSS CLKBUF_X1 
XU629 n608 n607 VDD VSS CLKBUF_X1 
XU630 n606 n608 VDD VSS INV_X32 
XU631 n607 n609 VDD VSS INV_X32 
XU632 c0_r4[9] n612 VDD VSS CLKBUF_X1 
XU633 n614 n613 VDD VSS CLKBUF_X1 
XU634 n612 n614 VDD VSS INV_X32 
XU635 n613 n615 VDD VSS INV_X32 
XU636 c0_r4[8] n616 VDD VSS CLKBUF_X1 
XU637 n618 n617 VDD VSS CLKBUF_X1 
XU638 n616 n618 VDD VSS INV_X32 
XU639 n617 n619 VDD VSS INV_X32 
XU640 c0_r4[7] n621 VDD VSS CLKBUF_X1 
XU641 n623 n622 VDD VSS CLKBUF_X1 
XU642 n621 n623 VDD VSS INV_X32 
XU643 n622 n624 VDD VSS INV_X32 
XU644 c0_r4[6] n625 VDD VSS CLKBUF_X1 
XU645 n627 n626 VDD VSS CLKBUF_X1 
XU646 n625 n627 VDD VSS INV_X32 
XU647 n626 n628 VDD VSS INV_X32 
XU648 c0_r4[5] n629 VDD VSS CLKBUF_X1 
XU649 n632 n631 VDD VSS CLKBUF_X1 
XU650 n629 n632 VDD VSS INV_X32 
XU651 n631 n633 VDD VSS INV_X32 
XU652 c0_r4[4] n634 VDD VSS CLKBUF_X1 
XU653 n636 n635 VDD VSS CLKBUF_X1 
XU654 n634 n636 VDD VSS INV_X32 
XU655 n635 n637 VDD VSS INV_X32 
XU656 c0_r4[3] n638 VDD VSS CLKBUF_X1 
XU657 n641 n639 VDD VSS CLKBUF_X1 
XU658 n638 n641 VDD VSS INV_X32 
XU659 n639 n642 VDD VSS INV_X32 
XU660 c0_r4[2] n643 VDD VSS CLKBUF_X1 
XU661 n645 n644 VDD VSS CLKBUF_X1 
XU662 n643 n645 VDD VSS INV_X32 
XU663 n644 n646 VDD VSS INV_X32 
XU664 c0_r4[1] n647 VDD VSS CLKBUF_X1 
XU665 n649 n648 VDD VSS CLKBUF_X1 
XU666 n647 n649 VDD VSS INV_X32 
XU667 n648 n651 VDD VSS INV_X32 
XU668 c0_r4[0] n652 VDD VSS CLKBUF_X1 
XU669 n654 n653 VDD VSS CLKBUF_X1 
XU670 n652 n654 VDD VSS INV_X32 
XU671 n653 n655 VDD VSS INV_X32 
XU672 sign_r[0] n656 VDD VSS CLKBUF_X1 
XU673 n658 n657 VDD VSS CLKBUF_X1 
XU674 n656 n658 VDD VSS INV_X32 
XU675 n657 n659 VDD VSS INV_X32 
XU676 sign_r[1] n661 VDD VSS CLKBUF_X1 
XU677 n663 n662 VDD VSS CLKBUF_X1 
XU678 n661 n663 VDD VSS INV_X32 
XU679 n662 n664 VDD VSS INV_X32 
XU680 sign_r[2] n665 VDD VSS CLKBUF_X1 
XU681 n667 n666 VDD VSS CLKBUF_X1 
XU682 n665 n667 VDD VSS INV_X32 
XU683 n666 n668 VDD VSS INV_X32 
XU684 sign_r[3] n669 VDD VSS CLKBUF_X1 
XU685 n672 n671 VDD VSS CLKBUF_X1 
XU686 n669 n672 VDD VSS INV_X32 
XU687 n671 n673 VDD VSS INV_X32 
XU688 sign_r[4] n674 VDD VSS CLKBUF_X1 
XU689 n676 n675 VDD VSS CLKBUF_X1 
XU690 n674 n676 VDD VSS INV_X32 
XU691 n675 n677 VDD VSS INV_X32 
XU692 n682 n678 VDD VSS BUF_X1 
XU693 n681 n679 VDD VSS CLKBUF_X1 
XU694 sign_r[5] n681 VDD VSS INV_X32 
XU695 n679 n682 VDD VSS INV_X32 
XU696 sign_r[6] n683 VDD VSS CLKBUF_X1 
XU697 n685 n684 VDD VSS CLKBUF_X1 
XU698 n683 n685 VDD VSS INV_X32 
XU699 n684 n686 VDD VSS INV_X32 
XU700 sign_r[7] n687 VDD VSS CLKBUF_X1 
XU701 n689 n688 VDD VSS CLKBUF_X1 
XU702 n687 n689 VDD VSS INV_X32 
XU703 n688 n691 VDD VSS INV_X32 
XU704 n695 n692 VDD VSS BUF_X1 
XU705 n694 n693 VDD VSS CLKBUF_X1 
XU706 N107 n694 VDD VSS INV_X32 
XU707 n693 n695 VDD VSS INV_X32 
XU708 N108 n696 VDD VSS CLKBUF_X1 
XU709 n698 n697 VDD VSS CLKBUF_X1 
XU710 n696 n698 VDD VSS INV_X32 
XU711 n697 n699 VDD VSS INV_X32 
XU712 valid_in_r[1] n701 VDD VSS CLKBUF_X1 
XU713 n703 n702 VDD VSS CLKBUF_X1 
XU714 n701 n703 VDD VSS INV_X32 
XU715 n702 n704 VDD VSS INV_X32 
XU716 N11010 n705 VDD VSS CLKBUF_X1 
XU717 n707 n706 VDD VSS CLKBUF_X1 
XU718 n705 n707 VDD VSS INV_X32 
XU719 n706 n708 VDD VSS INV_X32 
XU720 N111 n709 VDD VSS CLKBUF_X1 
XU721 n713 n712 VDD VSS CLKBUF_X1 
XU722 n709 n713 VDD VSS INV_X32 
XU723 n712 n714 VDD VSS INV_X32 
XU724 N112 n715 VDD VSS CLKBUF_X1 
XU725 n717 n716 VDD VSS CLKBUF_X1 
XU726 n715 n717 VDD VSS INV_X32 
XU727 n716 n718 VDD VSS INV_X32 
XU728 N113 n719 VDD VSS CLKBUF_X1 
XU729 n722 n721 VDD VSS CLKBUF_X1 
XU730 n719 n722 VDD VSS INV_X32 
XU731 n721 n723 VDD VSS INV_X32 
XU732 N114 n724 VDD VSS CLKBUF_X1 
XU733 n726 n725 VDD VSS CLKBUF_X1 
XU734 n724 n726 VDD VSS INV_X32 
XU735 n725 n727 VDD VSS INV_X32 
XU736 N115 n728 VDD VSS CLKBUF_X1 
XU737 n731 n729 VDD VSS CLKBUF_X1 
XU738 n728 n731 VDD VSS INV_X32 
XU739 n729 n732 VDD VSS INV_X32 
XU740 n736 n733 VDD VSS CLKBUF_X1 
XU741 n733 n734 VDD VSS INV_X32 
XU742 n734 n735 VDD VSS INV_X1 
XU743 n57 n736 VDD VSS INV_X1 
XU744 n735 n737 VDD VSS INV_X32 
XU745 n741 n738 VDD VSS CLKBUF_X1 
XU746 n742 n739 VDD VSS INV_X32 
XU747 n739 n741 VDD VSS INV_X1 
XU748 n28 n742 VDD VSS INV_X1 
XU749 n738 n743 VDD VSS INV_X32 
XU750 n746 n744 VDD VSS CLKBUF_X1 
XU751 n747 n745 VDD VSS INV_X32 
XU752 n745 n746 VDD VSS INV_X1 
XU753 n27 n747 VDD VSS INV_X1 
XU754 n744 n748 VDD VSS INV_X32 
XU755 n752 n749 VDD VSS CLKBUF_X1 
XU756 n753 n751 VDD VSS INV_X32 
XU757 n751 n752 VDD VSS INV_X1 
XU758 n26 n753 VDD VSS INV_X1 
XU759 n749 n754 VDD VSS INV_X32 
XU760 n759 n755 VDD VSS BUF_X1 
XU761 n758 n756 VDD VSS INV_X32 
XU762 n756 n757 VDD VSS INV_X1 
XU763 n25 n758 VDD VSS INV_X1 
XU764 n757 n759 VDD VSS INV_X32 
XU765 n764 n761 VDD VSS CLKBUF_X1 
XU766 n761 n762 VDD VSS INV_X32 
XU767 n762 n763 VDD VSS INV_X1 
XU768 n24 n764 VDD VSS INV_X1 
XU769 n763 n765 VDD VSS INV_X32 
XU770 n769 n766 VDD VSS CLKBUF_X1 
XU771 n766 n767 VDD VSS INV_X32 
XU772 n767 n768 VDD VSS INV_X1 
XU773 n23 n769 VDD VSS INV_X1 
XU774 n768 n771 VDD VSS INV_X32 
XU775 x_r2[7] n772 VDD VSS CLKBUF_X1 
XU776 n774 n773 VDD VSS CLKBUF_X1 
XU777 n772 n774 VDD VSS INV_X32 
XU778 n773 n775 VDD VSS INV_X32 
XU779 n777 n776 VDD VSS CLKBUF_X1 
XU780 n781 n777 VDD VSS INV_X1 
XU781 n776 n778 VDD VSS INV_X32 
XU782 N100 n779 VDD VSS INV_X1 
XU783 n779 n781 VDD VSS INV_X32 
XU784 x_r1[6] n782 VDD VSS CLKBUF_X1 
XU785 n784 n783 VDD VSS CLKBUF_X1 
XU786 n782 n784 VDD VSS INV_X32 
XU787 n783 n785 VDD VSS INV_X32 
XU788 x_r2[6] n786 VDD VSS CLKBUF_X1 
XU789 n788 n787 VDD VSS CLKBUF_X1 
XU790 n786 n788 VDD VSS INV_X32 
XU791 n787 n789 VDD VSS INV_X32 
XU792 n794 n791 VDD VSS CLKBUF_X1 
XU793 N101 n792 VDD VSS INV_X1 
XU794 n792 n793 VDD VSS INV_X32 
XU795 n793 n794 VDD VSS INV_X1 
XU796 n791 n795 VDD VSS INV_X32 
XU797 x_r1[5] n796 VDD VSS CLKBUF_X1 
XU798 n798 n797 VDD VSS CLKBUF_X1 
XU799 n796 n798 VDD VSS INV_X32 
XU800 n797 n799 VDD VSS INV_X32 
XU801 x_r2[5] n801 VDD VSS CLKBUF_X1 
XU802 n803 n802 VDD VSS CLKBUF_X1 
XU803 n801 n803 VDD VSS INV_X32 
XU804 n802 n804 VDD VSS INV_X32 
XU805 n806 n805 VDD VSS CLKBUF_X1 
XU806 N102 n806 VDD VSS INV_X1 
XU807 n805 n807 VDD VSS INV_X32 
XU808 n807 n808 VDD VSS INV_X1 
XU809 n808 n809 VDD VSS INV_X32 
XU810 x_r1[4] n812 VDD VSS CLKBUF_X1 
XU811 n814 n813 VDD VSS CLKBUF_X1 
XU812 n812 n814 VDD VSS INV_X32 
XU813 n813 n815 VDD VSS INV_X32 
XU814 x_r2[4] n816 VDD VSS CLKBUF_X1 
XU815 n818 n817 VDD VSS CLKBUF_X1 
XU816 n816 n818 VDD VSS INV_X32 
XU817 n817 n819 VDD VSS INV_X32 
XU818 n824 n821 VDD VSS CLKBUF_X1 
XU819 N103 n822 VDD VSS INV_X1 
XU820 n822 n823 VDD VSS INV_X32 
XU821 n823 n824 VDD VSS INV_X1 
XU822 n821 n825 VDD VSS INV_X32 
XU823 x_r1[3] n826 VDD VSS CLKBUF_X1 
XU824 n828 n827 VDD VSS CLKBUF_X1 
XU825 n826 n828 VDD VSS INV_X32 
XU826 n827 n829 VDD VSS INV_X32 
XU827 x_r2[3] n831 VDD VSS CLKBUF_X1 
XU828 n833 n832 VDD VSS CLKBUF_X1 
XU829 n831 n833 VDD VSS INV_X32 
XU830 n832 n834 VDD VSS INV_X32 
XU831 n837 n835 VDD VSS INV_X32 
XU832 n835 n836 VDD VSS INV_X1 
XU833 n841 n837 VDD VSS INV_X1 
XU834 n836 n838 VDD VSS INV_X32 
XU835 N104 n839 VDD VSS INV_X1 
XU836 n839 n841 VDD VSS INV_X32 
XU837 x_r1[2] n842 VDD VSS CLKBUF_X1 
XU838 n844 n843 VDD VSS CLKBUF_X1 
XU839 n842 n844 VDD VSS INV_X32 
XU840 n843 n845 VDD VSS INV_X32 
XU841 x_r2[2] n846 VDD VSS CLKBUF_X1 
XU842 n848 n847 VDD VSS CLKBUF_X1 
XU843 n846 n848 VDD VSS INV_X32 
XU844 n847 n849 VDD VSS INV_X32 
XU845 n854 n851 VDD VSS CLKBUF_X1 
XU846 N105 n852 VDD VSS INV_X1 
XU847 n852 n853 VDD VSS INV_X32 
XU848 n853 n854 VDD VSS INV_X1 
XU849 n851 n855 VDD VSS INV_X32 
XU850 x_r1[1] n856 VDD VSS CLKBUF_X1 
XU851 n858 n857 VDD VSS CLKBUF_X1 
XU852 n856 n858 VDD VSS INV_X32 
XU853 n857 n859 VDD VSS INV_X32 
XU854 x_r2[1] n861 VDD VSS CLKBUF_X1 
XU855 n863 n862 VDD VSS CLKBUF_X1 
XU856 n861 n863 VDD VSS INV_X32 
XU857 n862 n864 VDD VSS INV_X32 
XU858 n868 n865 VDD VSS INV_X1 
XU859 n865 n866 VDD VSS INV_X32 
XU860 n871 n867 VDD VSS INV_X1 
XU861 n867 n868 VDD VSS INV_X32 
XU862 N106 n869 VDD VSS INV_X1 
XU863 n869 n871 VDD VSS INV_X32 
XU864 x_r1[0] n872 VDD VSS CLKBUF_X1 
XU865 n874 n873 VDD VSS CLKBUF_X1 
XU866 n872 n874 VDD VSS INV_X32 
XU867 n873 n875 VDD VSS INV_X32 
XU868 x_r2[0] n876 VDD VSS CLKBUF_X1 
XU869 n878 n877 VDD VSS CLKBUF_X1 
XU870 n876 n878 VDD VSS INV_X32 
XU871 n877 n879 VDD VSS INV_X32 
XU872 x_r3[14] n881 VDD VSS CLKBUF_X1 
XU873 n883 n882 VDD VSS CLKBUF_X1 
XU874 n881 n883 VDD VSS INV_X32 
XU875 n882 n884 VDD VSS INV_X32 
XU876 x_r3[13] n885 VDD VSS CLKBUF_X1 
XU877 n887 n886 VDD VSS CLKBUF_X1 
XU878 n885 n887 VDD VSS INV_X32 
XU879 n886 n888 VDD VSS INV_X32 
XU880 x_r3[12] n889 VDD VSS CLKBUF_X1 
XU881 n892 n891 VDD VSS CLKBUF_X1 
XU882 n889 n892 VDD VSS INV_X32 
XU883 n891 n893 VDD VSS INV_X32 
XU884 x_r3[11] n894 VDD VSS CLKBUF_X1 
XU885 n896 n895 VDD VSS CLKBUF_X1 
XU886 n894 n896 VDD VSS INV_X32 
XU887 n895 n897 VDD VSS INV_X32 
XU888 x_r3[10] n898 VDD VSS CLKBUF_X1 
XU889 n901 n899 VDD VSS CLKBUF_X1 
XU890 n898 n901 VDD VSS INV_X32 
XU891 n899 n902 VDD VSS INV_X32 
XU892 x_r3[9] n903 VDD VSS CLKBUF_X1 
XU893 n905 n904 VDD VSS CLKBUF_X1 
XU894 n903 n905 VDD VSS INV_X32 
XU895 n904 n906 VDD VSS INV_X32 
XU896 x_r3[8] n907 VDD VSS CLKBUF_X1 
XU897 n909 n908 VDD VSS CLKBUF_X1 
XU898 n907 n909 VDD VSS INV_X32 
XU899 n908 n912 VDD VSS INV_X32 
XU900 x_r3[7] n913 VDD VSS CLKBUF_X1 
XU901 n915 n914 VDD VSS CLKBUF_X1 
XU902 n913 n915 VDD VSS INV_X32 
XU903 n914 n916 VDD VSS INV_X32 
XU904 x_r3[6] n917 VDD VSS CLKBUF_X1 
XU905 n919 n918 VDD VSS CLKBUF_X1 
XU906 n917 n919 VDD VSS INV_X32 
XU907 n918 n921 VDD VSS INV_X32 
XU908 x_r3[5] n922 VDD VSS CLKBUF_X1 
XU909 n924 n923 VDD VSS CLKBUF_X1 
XU910 n922 n924 VDD VSS INV_X32 
XU911 n923 n925 VDD VSS INV_X32 
XU912 x_r3[4] n926 VDD VSS CLKBUF_X1 
XU913 n928 n927 VDD VSS CLKBUF_X1 
XU914 n926 n928 VDD VSS INV_X32 
XU915 n927 n929 VDD VSS INV_X32 
XU916 x_r3[3] n931 VDD VSS CLKBUF_X1 
XU917 n933 n932 VDD VSS CLKBUF_X1 
XU918 n931 n933 VDD VSS INV_X32 
XU919 n932 n934 VDD VSS INV_X32 
XU920 x_r3[2] n935 VDD VSS CLKBUF_X1 
XU921 n937 n936 VDD VSS CLKBUF_X1 
XU922 n935 n937 VDD VSS INV_X32 
XU923 n936 n938 VDD VSS INV_X32 
XU924 x_r3[1] n939 VDD VSS CLKBUF_X1 
XU925 n942 n941 VDD VSS CLKBUF_X1 
XU926 n939 n942 VDD VSS INV_X32 
XU927 n941 n943 VDD VSS INV_X32 
XU928 x_r3[0] n944 VDD VSS CLKBUF_X1 
XU929 n946 n945 VDD VSS CLKBUF_X1 
XU930 n944 n946 VDD VSS INV_X32 
XU931 n945 n947 VDD VSS INV_X32 
XU932 c0_r1[17] n948 VDD VSS CLKBUF_X1 
XU933 n951 n949 VDD VSS CLKBUF_X1 
XU934 n948 n951 VDD VSS INV_X32 
XU935 n949 n952 VDD VSS INV_X32 
XU936 c0_r2[17] n953 VDD VSS CLKBUF_X1 
XU937 n955 n954 VDD VSS CLKBUF_X1 
XU938 n953 n955 VDD VSS INV_X32 
XU939 n954 n956 VDD VSS INV_X32 
XU940 c0_r3[17] n957 VDD VSS CLKBUF_X1 
XU941 n959 n958 VDD VSS CLKBUF_X1 
XU942 n957 n959 VDD VSS INV_X32 
XU943 n958 n960 VDD VSS INV_X32 
XU944 c0_r1[16] n961 VDD VSS CLKBUF_X1 
XU945 n963 n962 VDD VSS CLKBUF_X1 
XU946 n961 n963 VDD VSS INV_X32 
XU947 n962 n964 VDD VSS INV_X32 
XU948 c0_r2[16] n965 VDD VSS CLKBUF_X1 
XU949 n967 n966 VDD VSS CLKBUF_X1 
XU950 n965 n967 VDD VSS INV_X32 
XU951 n966 n968 VDD VSS INV_X32 
XU952 c0_r3[16] n969 VDD VSS CLKBUF_X1 
XU953 n971 n970 VDD VSS CLKBUF_X1 
XU954 n969 n971 VDD VSS INV_X32 
XU955 n970 n972 VDD VSS INV_X32 
XU956 c0_r1[15] n973 VDD VSS CLKBUF_X1 
XU957 n975 n974 VDD VSS CLKBUF_X1 
XU958 n973 n975 VDD VSS INV_X32 
XU959 n974 n976 VDD VSS INV_X32 
XU960 c0_r2[15] n977 VDD VSS CLKBUF_X1 
XU961 n979 n978 VDD VSS CLKBUF_X1 
XU962 n977 n979 VDD VSS INV_X32 
XU963 n978 n981 VDD VSS INV_X32 
XU964 c0_r3[15] n982 VDD VSS CLKBUF_X1 
XU965 n984 n983 VDD VSS CLKBUF_X1 
XU966 n982 n984 VDD VSS INV_X32 
XU967 n983 n985 VDD VSS INV_X32 
XU968 c0_r1[14] n986 VDD VSS CLKBUF_X1 
XU969 n988 n987 VDD VSS CLKBUF_X1 
XU970 n986 n988 VDD VSS INV_X32 
XU971 n987 n989 VDD VSS INV_X32 
XU972 c0_r2[14] n991 VDD VSS CLKBUF_X1 
XU973 n993 n992 VDD VSS CLKBUF_X1 
XU974 n991 n993 VDD VSS INV_X32 
XU975 n992 n994 VDD VSS INV_X32 
XU976 c0_r3[14] n995 VDD VSS CLKBUF_X1 
XU977 n997 n996 VDD VSS CLKBUF_X1 
XU978 n995 n997 VDD VSS INV_X32 
XU979 n996 n998 VDD VSS INV_X32 
XU980 c0_r1[13] n999 VDD VSS CLKBUF_X1 
XU981 n1002 n1001 VDD VSS CLKBUF_X1 
XU982 n999 n1002 VDD VSS INV_X32 
XU983 n1001 n1003 VDD VSS INV_X32 
XU984 c0_r2[13] n1004 VDD VSS CLKBUF_X1 
XU985 n1006 n1005 VDD VSS CLKBUF_X1 
XU986 n1004 n1006 VDD VSS INV_X32 
XU987 n1005 n1007 VDD VSS INV_X32 
XU988 c0_r3[13] n1008 VDD VSS CLKBUF_X1 
XU989 n1012 n1009 VDD VSS CLKBUF_X1 
XU990 n1008 n1012 VDD VSS INV_X32 
XU991 n1009 n1013 VDD VSS INV_X32 
XU992 c0_r1[12] n1014 VDD VSS CLKBUF_X1 
XU993 n1016 n1015 VDD VSS CLKBUF_X1 
XU994 n1014 n1016 VDD VSS INV_X32 
XU995 n1015 n1017 VDD VSS INV_X32 
XU996 c0_r2[12] n1018 VDD VSS CLKBUF_X1 
XU997 n1021 n1019 VDD VSS CLKBUF_X1 
XU998 n1018 n1021 VDD VSS INV_X32 
XU999 n1019 n1022 VDD VSS INV_X32 
XU1000 c0_r3[12] n1023 VDD VSS CLKBUF_X1 
XU1001 n1025 n1024 VDD VSS CLKBUF_X1 
XU1002 n1023 n1025 VDD VSS INV_X32 
XU1003 n1024 n1026 VDD VSS INV_X32 
XU1004 c0_r1[11] n1027 VDD VSS CLKBUF_X1 
XU1005 n1029 n1028 VDD VSS CLKBUF_X1 
XU1006 n1027 n1029 VDD VSS INV_X32 
XU1007 n1028 n1031 VDD VSS INV_X32 
XU1008 c0_r2[11] n1032 VDD VSS CLKBUF_X1 
XU1009 n1034 n1033 VDD VSS CLKBUF_X1 
XU1010 n1032 n1034 VDD VSS INV_X32 
XU1011 n1033 n1035 VDD VSS INV_X32 
XU1012 c0_r3[11] n1036 VDD VSS CLKBUF_X1 
XU1013 n1038 n1037 VDD VSS CLKBUF_X1 
XU1014 n1036 n1038 VDD VSS INV_X32 
XU1015 n1037 n1039 VDD VSS INV_X32 
XU1016 c0_r1[10] n1041 VDD VSS CLKBUF_X1 
XU1017 n1043 n1042 VDD VSS CLKBUF_X1 
XU1018 n1041 n1043 VDD VSS INV_X32 
XU1019 n1042 n1044 VDD VSS INV_X32 
XU1020 c0_r2[10] n1045 VDD VSS CLKBUF_X1 
XU1021 n1047 n1046 VDD VSS CLKBUF_X1 
XU1022 n1045 n1047 VDD VSS INV_X32 
XU1023 n1046 n1048 VDD VSS INV_X32 
XU1024 n1053 n1049 VDD VSS BUF_X1 
XU1025 n1052 n1051 VDD VSS CLKBUF_X1 
XU1026 c0_r3[10] n1052 VDD VSS INV_X32 
XU1027 n1051 n1053 VDD VSS INV_X32 
XU1028 c0_r1[9] n1054 VDD VSS CLKBUF_X1 
XU1029 n1900 n1055 VDD VSS CLKBUF_X1 
XU1030 n1054 n1056 VDD VSS INV_X32 
XU1031 n1055 n1057 VDD VSS INV_X32 
XU1032 c0_r2[9] n1058 VDD VSS CLKBUF_X1 
XU1033 n1061 n1059 VDD VSS CLKBUF_X1 
XU1034 n1058 n1061 VDD VSS INV_X32 
XU1035 n1059 n1062 VDD VSS INV_X32 
XU1036 c0_r3[9] n1063 VDD VSS CLKBUF_X1 
XU1037 n1065 n1064 VDD VSS CLKBUF_X1 
XU1038 n1063 n1065 VDD VSS INV_X32 
XU1039 n1064 n1066 VDD VSS INV_X32 
XU1040 c0_r1[8] n1067 VDD VSS CLKBUF_X1 
XU1041 n1069 n1068 VDD VSS CLKBUF_X1 
XU1042 n1067 n1069 VDD VSS INV_X32 
XU1043 n1068 n1071 VDD VSS INV_X32 
XU1044 N11000 n1072 VDD VSS INV_X1 
XU1045 n1072 n1073 VDD VSS INV_X32 
XU1046 n1077 n1074 VDD VSS INV_X1 
XU1047 n1074 n1075 VDD VSS INV_X32 
XU1048 N10 n1076 VDD VSS INV_X1 
XU1049 n1076 n1077 VDD VSS INV_X32 
XU1050 N900 n1078 VDD VSS INV_X1 
XU1051 n1078 n1079 VDD VSS INV_X32 
XU1052 N8 n1081 VDD VSS BUF_X1 
XU1053 N700 n1082 VDD VSS CLKBUF_X1 
XU1054 N74 n1083 VDD VSS CLKBUF_X1 
XU1055 n1117 n1084 VDD VSS BUF_X1 
XU1056 N7010 n1085 VDD VSS BUF_X1 
XU1057 n7210 n1086 VDD VSS BUF_X1 
XU1058 num_lzd_r[3] n1087 VDD VSS INV_X1 
XU1059 n1087 n1088 VDD VSS INV_X32 
XU1060 n1010 n1089 VDD VSS INV_X1 
XU1061 n1089 n1091 VDD VSS INV_X32 
XU1062 n205 n10921 VDD VSS CLKBUF_X1 
XU1063 n810 n1093 VDD VSS CLKBUF_X1 
XU1064 n1110 n1094 VDD VSS INV_X1 
XU1065 n1094 n1095 VDD VSS INV_X16 
XU1066 n143 n1096 VDD VSS CLKBUF_X1 
XU1067 num_lzd_r[5] n1097 VDD VSS INV_X1 
XU1068 n1097 n1098 VDD VSS INV_X32 
XU1069 num_lzd_r[4] n1099 VDD VSS INV_X32 
XU1070 n1099 n1101 VDD VSS INV_X1 
XU1071 N65 n1102 VDD VSS INV_X1 
XU1072 n46 n1104 VDD VSS INV_X1 
XU1073 n1104 n1105 VDD VSS INV_X32 
XU1074 n1105 n1106 VDD VSS INV_X1 
XU1075 n1106 n1107 VDD VSS INV_X32 
XU1076 N64 n1108 VDD VSS INV_X1 
XU1077 n48 n1112 VDD VSS INV_X1 
XU1078 n1112 n1113 VDD VSS INV_X32 
XU1079 n1113 n1114 VDD VSS INV_X1 
XU1080 n1114 n1115 VDD VSS INV_X32 
XU1081 n50 n1116 VDD VSS INV_X32 
XU1082 n1122 n1118 VDD VSS INV_X1 
XU1083 n1118 n1119 VDD VSS INV_X32 
XU1084 n49 n1121 VDD VSS INV_X1 
XU1085 n1121 n1122 VDD VSS INV_X32 
XU1086 n1126 n1123 VDD VSS CLKBUF_X1 
XU1087 n910 n1124 VDD VSS INV_X1 
XU1088 n1124 n1125 VDD VSS INV_X32 
XU1089 n1093 n1126 VDD VSS INV_X32 
XU1090 N611 n1128 VDD VSS INV_X1 
XU1091 n1128 n1129 VDD VSS INV_X16 
XU1092 n53 n1130 VDD VSS INV_X1 
XU1093 n1130 n1131 VDD VSS INV_X32 
XU1094 n1131 n1132 VDD VSS INV_X1 
XU1095 n1132 n1133 VDD VSS INV_X32 
XU1096 n1137 n1134 VDD VSS BUF_X1 
XU1097 n1136 n1135 VDD VSS CLKBUF_X1 
XU1098 N600 n1136 VDD VSS INV_X32 
XU1099 n1135 n1137 VDD VSS INV_X32 
XU1100 N76 n1138 VDD VSS CLKBUF_X1 
XU1101 n1140 n1139 VDD VSS CLKBUF_X1 
XU1102 n1138 n1140 VDD VSS INV_X32 
XU1103 n1139 n1141 VDD VSS INV_X32 
XU1104 n1145 n1142 VDD VSS BUF_X1 
XU1105 n1144 n1143 VDD VSS CLKBUF_X1 
XU1106 N75 n1144 VDD VSS INV_X32 
XU1107 n1143 n1145 VDD VSS INV_X32 
XU1108 N91 n1146 VDD VSS CLKBUF_X1 
XU1109 n1148 n1147 VDD VSS CLKBUF_X1 
XU1110 n1146 n1148 VDD VSS INV_X32 
XU1111 n1147 n1149 VDD VSS INV_X32 
XU1112 N9010 n1150 VDD VSS CLKBUF_X1 
XU1113 n1152 n1151 VDD VSS CLKBUF_X1 
XU1114 n1150 n1152 VDD VSS INV_X32 
XU1115 n1151 n1153 VDD VSS INV_X32 
XU1116 N89 n1154 VDD VSS CLKBUF_X1 
XU1117 n1156 n1155 VDD VSS CLKBUF_X1 
XU1118 n1154 n1156 VDD VSS INV_X32 
XU1119 n1155 n1157 VDD VSS INV_X32 
XU1120 N88 n1158 VDD VSS INV_X1 
XU1121 n1930 n1159 VDD VSS INV_X32 
XU1122 N87 n1160 VDD VSS CLKBUF_X1 
XU1123 n1162 n1161 VDD VSS CLKBUF_X1 
XU1124 n1160 n1162 VDD VSS INV_X32 
XU1125 n1161 n1163 VDD VSS INV_X32 
XU1126 n1165 n1164 VDD VSS CLKBUF_X1 
XU1127 N86 n1165 VDD VSS INV_X32 
XU1128 n1164 n1166 VDD VSS INV_X32 
XU1129 n1170 n1167 VDD VSS CLKBUF_X1 
XU1130 n1169 n1168 VDD VSS CLKBUF_X1 
XU1131 N85 n1169 VDD VSS INV_X32 
XU1132 n1168 n1170 VDD VSS INV_X32 
XU1133 N84 n1171 VDD VSS CLKBUF_X1 
XU1134 n1173 n1172 VDD VSS CLKBUF_X1 
XU1135 n1171 n1173 VDD VSS INV_X32 
XU1136 n1172 n1174 VDD VSS INV_X32 
XU1137 N83 n1175 VDD VSS CLKBUF_X1 
XU1138 n1177 n1176 VDD VSS CLKBUF_X1 
XU1139 n1175 n1177 VDD VSS INV_X32 
XU1140 n1176 n1178 VDD VSS INV_X32 
XU1141 N82 n1179 VDD VSS CLKBUF_X1 
XU1142 n1181 n1180 VDD VSS CLKBUF_X1 
XU1143 n1179 n1181 VDD VSS INV_X32 
XU1144 n1180 n1182 VDD VSS INV_X32 
XU1145 N81 n1183 VDD VSS CLKBUF_X1 
XU1146 n1185 n1184 VDD VSS CLKBUF_X1 
XU1147 n1183 n1185 VDD VSS INV_X32 
XU1148 n1184 n1186 VDD VSS INV_X32 
XU1149 N79 n1187 VDD VSS CLKBUF_X1 
XU1150 n1189 n1188 VDD VSS CLKBUF_X1 
XU1151 n1187 n1189 VDD VSS INV_X32 
XU1152 n1188 n1190 VDD VSS INV_X32 
XU1153 n1194 n1191 VDD VSS BUF_X1 
XU1154 n1193 n1192 VDD VSS CLKBUF_X1 
XU1155 N78 n1193 VDD VSS INV_X32 
XU1156 n1192 n1194 VDD VSS INV_X32 
XU1157 n1198 n1195 VDD VSS BUF_X1 
XU1158 n1197 n1196 VDD VSS CLKBUF_X1 
XU1159 N77 n1197 VDD VSS INV_X32 
XU1160 n1196 n1198 VDD VSS INV_X32 
XU1161 n1201 n1199 VDD VSS INV_X32 
XU1162 n1199 n1200 VDD VSS INV_X1 
XU1163 n1204 n1201 VDD VSS INV_X1 
XU1164 n1200 n1202 VDD VSS INV_X32 
XU1165 N92 n1203 VDD VSS INV_X1 
XU1166 n1203 n1204 VDD VSS INV_X32 
XU1167 x_r1[14] n1205 VDD VSS CLKBUF_X1 
XU1168 n1207 n1206 VDD VSS CLKBUF_X1 
XU1169 n1205 n1207 VDD VSS INV_X32 
XU1170 n1206 n1208 VDD VSS INV_X32 
XU1171 x_r2[14] n1209 VDD VSS CLKBUF_X1 
XU1172 n1211 n1210 VDD VSS CLKBUF_X1 
XU1173 n1209 n1211 VDD VSS INV_X32 
XU1174 n1210 n1212 VDD VSS INV_X32 
XU1175 n1215 n1213 VDD VSS INV_X32 
XU1176 n1213 n1214 VDD VSS INV_X1 
XU1177 n1218 n1215 VDD VSS INV_X1 
XU1178 n1214 n1216 VDD VSS INV_X32 
XU1179 N93 n1217 VDD VSS INV_X1 
XU1180 n1217 n1218 VDD VSS INV_X32 
XU1181 x_r1[13] n1219 VDD VSS CLKBUF_X1 
XU1182 n1221 n1220 VDD VSS CLKBUF_X1 
XU1183 n1219 n1221 VDD VSS INV_X32 
XU1184 n1220 n1222 VDD VSS INV_X32 
XU1185 x_r2[13] n1223 VDD VSS CLKBUF_X1 
XU1186 n1225 n1224 VDD VSS CLKBUF_X1 
XU1187 n1223 n1225 VDD VSS INV_X32 
XU1188 n1224 n1226 VDD VSS INV_X32 
XU1189 n1228 n1227 VDD VSS CLKBUF_X1 
XU1190 n1231 n1228 VDD VSS INV_X1 
XU1191 n1227 n1229 VDD VSS INV_X32 
XU1192 N94 n1230 VDD VSS INV_X1 
XU1193 n1230 n1231 VDD VSS INV_X32 
XU1194 x_r1[12] n1232 VDD VSS CLKBUF_X1 
XU1195 n1234 n1233 VDD VSS CLKBUF_X1 
XU1196 n1232 n1234 VDD VSS INV_X32 
XU1197 n1233 n1235 VDD VSS INV_X32 
XU1198 x_r2[12] n1236 VDD VSS CLKBUF_X1 
XU1199 n1238 n1237 VDD VSS CLKBUF_X1 
XU1200 n1236 n1238 VDD VSS INV_X32 
XU1201 n1237 n1239 VDD VSS INV_X32 
XU1202 n1242 n1240 VDD VSS INV_X32 
XU1203 n1240 n1241 VDD VSS INV_X1 
XU1204 N95 n1242 VDD VSS INV_X1 
XU1205 n1241 n1243 VDD VSS INV_X32 
XU1206 n1243 n1244 VDD VSS INV_X1 
XU1207 n1244 n1245 VDD VSS INV_X32 
XU1208 x_r1[11] n1246 VDD VSS CLKBUF_X1 
XU1209 n1248 n1247 VDD VSS CLKBUF_X1 
XU1210 n1246 n1248 VDD VSS INV_X32 
XU1211 n1247 n1249 VDD VSS INV_X32 
XU1212 x_r2[11] n1250 VDD VSS CLKBUF_X1 
XU1213 n1252 n1251 VDD VSS CLKBUF_X1 
XU1214 n1250 n1252 VDD VSS INV_X32 
XU1215 n1251 n1253 VDD VSS INV_X32 
XU1216 n1255 n1254 VDD VSS CLKBUF_X1 
XU1217 N96 n1255 VDD VSS INV_X1 
XU1218 n1254 n1256 VDD VSS INV_X32 
XU1219 n1256 n1257 VDD VSS INV_X1 
XU1220 n1257 n1258 VDD VSS INV_X32 
XU1221 x_r1[10] n1259 VDD VSS CLKBUF_X1 
XU1222 n1261 n1260 VDD VSS CLKBUF_X1 
XU1223 n1259 n1261 VDD VSS INV_X32 
XU1224 n1260 n1262 VDD VSS INV_X32 
XU1225 x_r2[10] n1263 VDD VSS CLKBUF_X1 
XU1226 n1265 n1264 VDD VSS CLKBUF_X1 
XU1227 n1263 n1265 VDD VSS INV_X32 
XU1228 n1264 n1266 VDD VSS INV_X32 
XU1229 n1270 n1267 VDD VSS INV_X1 
XU1231 n1272 n1269 VDD VSS INV_X1 
XU1232 n1269 n1270 VDD VSS INV_X32 
XU1233 N97 n1271 VDD VSS INV_X1 
XU1234 n1271 n1272 VDD VSS INV_X32 
XU1235 x_r1[9] n1273 VDD VSS CLKBUF_X1 
XU1236 n1275 n1274 VDD VSS CLKBUF_X1 
XU1237 n1273 n1275 VDD VSS INV_X32 
XU1238 n1274 n1276 VDD VSS INV_X32 
XU1239 x_r2[9] n1277 VDD VSS CLKBUF_X1 
XU1240 n1279 n1278 VDD VSS CLKBUF_X1 
XU1241 n1277 n1279 VDD VSS INV_X32 
XU1242 n1278 n1280 VDD VSS INV_X32 
XU1243 n1284 n1281 VDD VSS CLKBUF_X1 
XU1244 N98 n1282 VDD VSS INV_X1 
XU1245 n1282 n1283 VDD VSS INV_X32 
XU1246 n1283 n1284 VDD VSS INV_X1 
XU1247 n1281 n1285 VDD VSS INV_X32 
XU1248 x_r1[8] n1286 VDD VSS CLKBUF_X1 
XU1249 n1288 n1287 VDD VSS CLKBUF_X1 
XU1250 n1286 n1288 VDD VSS INV_X32 
XU1251 n1287 n1289 VDD VSS INV_X32 
XU1252 x_r2[8] n1290 VDD VSS CLKBUF_X1 
XU1253 n1292 n1291 VDD VSS CLKBUF_X1 
XU1254 n1290 n1292 VDD VSS INV_X32 
XU1255 n1291 n1293 VDD VSS INV_X32 
XU1256 n1298 n1294 VDD VSS INV_X32 
XU1257 n1294 n1295 VDD VSS INV_X1 
XU1258 N99 n1296 VDD VSS INV_X1 
XU1259 n1296 n1297 VDD VSS INV_X32 
XU1260 n1297 n1298 VDD VSS INV_X1 
XU1261 n1295 n1299 VDD VSS INV_X32 
XU1262 x_r1[7] n1300 VDD VSS CLKBUF_X1 
XU1263 n1302 n1301 VDD VSS CLKBUF_X1 
XU1264 n1300 n1302 VDD VSS INV_X32 
XU1265 n1301 n1303 VDD VSS INV_X32 
XU1230 n1267 n1268 VDD VSS INV_X16 
XU1266 n446 n1304 VDD VSS BUF_X1 
XU1267 N127 n1305 VDD VSS BUF_X1 
XU1268 n1268 n1306 VDD VSS BUF_X1 
XU1269 n1306 n1307 VDD VSS BUF_X1 
XU1294 n135 n1332 VDD VSS BUF_X1 
XU1295 n425 n1333 VDD VSS BUF_X1 
XU1296 n1285 n1334 VDD VSS BUF_X1 
XU1270 N121 n1335 VDD VSS BUF_X1 
XU1271 n1335 n1336 VDD VSS BUF_X1 
Xu_gng_lzd num_lzd[5] num_lzd[4] num_lzd[3] num_lzd[2] num_lzd[1] num_lzd[0] VDD 
+ VSS data_in[63] data_in[62] data_in[61] data_in[60] data_in[59] data_in[58] data_in[57] 
+ data_in[56] data_in[55] data_in[54] data_in[53] data_in[52] data_in[51] data_in[50] 
+ data_in[49] data_in[48] data_in[47] data_in[46] data_in[45] data_in[44] data_in[43] 
+ data_in[42] data_in[41] data_in[40] data_in[39] data_in[38] data_in[37] data_in[36] 
+ data_in[35] data_in[34] data_in[33] data_in[32] data_in[31] data_in[30] data_in[29] 
+ data_in[28] data_in[27] data_in[26] data_in[25] data_in[24] data_in[23] data_in[22] 
+ data_in[21] data_in[20] data_in[19] data_in[18] data_in[17] data_in[16] data_in[15] 
+ data_in[14] data_in[13] data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] 
+ data_in[7] data_in[6] data_in[5] data_in[4] data_in[3] gng_lzd 
Xu_gng_coef c2[16] c2[15] c2[14] c2[13] c2[12] c2[11] c2[10] c2[9] c2[8] c2[7] c2[6] 
+ c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] n6310 VDD VSS c1[17] c1[16] c1[15] c1[14] 
+ c1[13] c1[12] c1[11] c1[10] c1[9] c1[8] c1[7] c1[6] c1[5] c1[4] c1[3] c1[2] c1[1] 
+ c1[0] c0[17] c0[16] c0[15] c0[14] c0[13] c0[12] c0[11] c0[10] c0[9] c0[8] c0[7] 
+ c0[6] c0[5] c0[4] c0[3] c0[2] c0[1] c0[0] n6810 n10921 n7011 n1096 n7210 n7310 
+ n202 n207 n132 n133 n143 n142 n205 n1332 n63_G2B1I8 n63_G2B1I2 gng_coef 
Xu_gng_smul_16_18_sadd_37 sum1[37] sum1[36] sum1[35] sum1[34] sum1[33] sum1[32] 
+ sum1[31] sum1[30] sum1[29] sum1[28] sum1[27] sum1[26] sum1[25] sum1[24] sum1[23] 
+ sum1[22] sum1[21] sum1[20] SYNOPSYS_UNCONNECTED_26 SYNOPSYS_UNCONNECTED_25 SYNOPSYS_UNCONNECTED_24 
+ SYNOPSYS_UNCONNECTED_34 SYNOPSYS_UNCONNECTED_33 SYNOPSYS_UNCONNECTED_32 SYNOPSYS_UNCONNECTED_31 
+ SYNOPSYS_UNCONNECTED_30 SYNOPSYS_UNCONNECTED_29 SYNOPSYS_UNCONNECTED_28 SYNOPSYS_UNCONNECTED_27 
+ SYNOPSYS_UNCONNECTED_42 SYNOPSYS_UNCONNECTED_41 SYNOPSYS_UNCONNECTED_40 SYNOPSYS_UNCONNECTED_39 
+ SYNOPSYS_UNCONNECTED_38 SYNOPSYS_UNCONNECTED_37 SYNOPSYS_UNCONNECTED_36 SYNOPSYS_UNCONNECTED_35 
+ SYNOPSYS_UNCONNECTED_43 n10920 VDD VSS n214 n218 n222 n226 n230 n234 n145 n242 
+ n246 n250 n1470 n258 n262 n266 n270 n148 n278 n282 VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS c2[16] c2[15] c2[14] c2[13] 
+ c2[12] c2[11] c2[10] c2[9] c2[8] c2[7] c2[6] c2[5] c2[4] c2[3] c2[2] c2[1] c2[0] 
+ VSS n1208 n1222 n1235 n1249 n1262 n1276 n209 n1303 n785 n210 n815 n829 n845 n859 
+ n875 gng_smul_16_18_sadd_37 
Xu_gng_smul_16_18 SYNOPSYS_UNCONNECTED_4 mul1[32] mul1[31] mul1[30] mul1[29] mul1[28] 
+ mul1[27] mul1[26] mul1[25] mul1[24] mul1[23] mul1[22] mul1[21] mul1[20] mul1[19] 
+ SYNOPSYS_UNCONNECTED_9 SYNOPSYS_UNCONNECTED_8 SYNOPSYS_UNCONNECTED_7 SYNOPSYS_UNCONNECTED_6 
+ SYNOPSYS_UNCONNECTED_5 SYNOPSYS_UNCONNECTED_17 SYNOPSYS_UNCONNECTED_16 SYNOPSYS_UNCONNECTED_15 
+ SYNOPSYS_UNCONNECTED_14 SYNOPSYS_UNCONNECTED_13 SYNOPSYS_UNCONNECTED_12 SYNOPSYS_UNCONNECTED_11 
+ SYNOPSYS_UNCONNECTED_10 SYNOPSYS_UNCONNECTED_23 SYNOPSYS_UNCONNECTED_22 SYNOPSYS_UNCONNECTED_21 
+ SYNOPSYS_UNCONNECTED_20 SYNOPSYS_UNCONNECTED_19 SYNOPSYS_UNCONNECTED_18 n6111 
+ VDD VSS sum1[37] sum1[36] sum1[35] sum1[34] sum1[33] sum1[32] sum1[31] sum1[30] 
+ sum1[29] sum1[28] sum1[27] sum1[26] sum1[25] sum1[24] sum1[23] sum1[22] sum1[21] 
+ sum1[20] VSS n286 n290 n294 n298 n302 n306 n310 n314 n318 n322 n326 n330 n334 
+ n338 n342 gng_smul_16_18 
Xadd_219 N1810 N1800 N1790 N1780 N1770 N1760 N1750 N1740 N1730 N1720 N1710 N1700 
+ N1690 N1680 N1670 SYNOPSYS_UNCONNECTED_3 VDD n29 n30 n31 n32 n33 n34 n35 n36 n37 
+ n38 n39 n40 n41 n42 n43 VDD VSS gng_interp_DW01_inc_0 
Xadd_199 N131 N130 N129 N128 N127 N126 N125 N124 N123 N122 N121 N120 N119 N118 N117 
+ N116 SYNOPSYS_UNCONNECTED_2 SYNOPSYS_UNCONNECTED_1 VSS SYNOPSYS_UNCONNECTED_273 
+ mul1[32] mul1[32] mul1[32] mul1[32] mul1[32] mul1[31] mul1[30] mul1[29] mul1[28] 
+ mul1[27] mul1[26] mul1[25] mul1[24] mul1[23] mul1[22] mul1[21] mul1[20] mul1[19] 
+ c0_r5[17] c0_r5[16] c0_r5[15] c0_r5[14] c0_r5[13] c0_r5[12] c0_r5[11] c0_r5[10] 
+ c0_r5[9] c0_r5[8] c0_r5[7] c0_r5[6] c0_r5[5] c0_r5[4] c0_r5[3] c0_r5[2] c0_r5[1] 
+ c0_r5[0] VDD VSS gng_interp_DW01_add_1 
.ENDS

.SUBCKT gng data_out[15] data_out[14] data_out[13] data_out[12] data_out[11] data_out[10] 
+ data_out[9] data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] data_out[3] 
+ data_out[2] data_out[1] data_out[0] valid_out ce rstn clk 
Xxofiller_FILLCELL_X2_8943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1099 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1098 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1097 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1096 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1095 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1094 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1093 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1092 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1091 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1090 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1089 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1088 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1087 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1086 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1085 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1084 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1083 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1082 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1081 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1080 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1079 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1078 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1077 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1076 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1075 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1074 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1073 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1072 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1071 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1070 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1069 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1068 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1067 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1066 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1065 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1064 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1063 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1062 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1061 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1060 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1059 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1058 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1057 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1056 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1055 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1054 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1053 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1052 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1051 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1050 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1049 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1048 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1047 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1046 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1045 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1044 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1043 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1042 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1041 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1040 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1039 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1038 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1037 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1036 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1035 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1034 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1033 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1032 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1031 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1030 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1029 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1028 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1027 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1026 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1025 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1024 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1023 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1022 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1021 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1020 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1019 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1018 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1017 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1016 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1015 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1014 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1013 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1012 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1011 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1010 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1009 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1008 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1007 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1006 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1005 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1004 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1003 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1002 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1001 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1000 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_999 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_998 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_997 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_996 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_995 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_994 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_993 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_992 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_991 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_990 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_989 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_988 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_987 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_986 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_985 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_984 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_983 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_982 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_981 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_980 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_979 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_978 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_977 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_976 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_975 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_974 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_973 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_972 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_971 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_970 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_969 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_968 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_967 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_966 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_965 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_964 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_963 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_962 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_961 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_960 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_959 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_958 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_957 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_956 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_955 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_954 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_953 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_952 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_951 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_950 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_949 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_948 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_947 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_946 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_945 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_944 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_943 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_942 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_941 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_940 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_939 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_938 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_937 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_936 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_935 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_934 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_933 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_932 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_931 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_930 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_929 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_928 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_927 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_926 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_925 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_924 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_923 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_922 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_921 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_920 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_919 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_918 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_917 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_916 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_915 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_914 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_913 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_912 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_911 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_910 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_909 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_908 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_907 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_906 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_905 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_904 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_903 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_902 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_901 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_900 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_899 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_898 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_897 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_896 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_895 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_894 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_893 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_892 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_891 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_890 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_889 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_888 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_887 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_886 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_885 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_884 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_883 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_882 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_881 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_880 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_879 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_878 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_877 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_876 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_875 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_874 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_873 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_872 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_871 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_870 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_869 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_868 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_867 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_866 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_865 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_864 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_863 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_862 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_861 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_860 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_859 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_858 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_857 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_856 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_855 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_854 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_853 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_852 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_851 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_850 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_849 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_848 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_847 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_846 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_845 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_844 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_843 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_842 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_841 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_840 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_839 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_838 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_837 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_836 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_835 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_834 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_833 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_832 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_831 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_830 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_829 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_828 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_827 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_826 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_825 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_824 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_823 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_822 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_821 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_820 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_819 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_818 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_817 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_816 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_815 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_814 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_813 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_812 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_811 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_810 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_809 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_808 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_807 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_806 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_805 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_804 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_803 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_802 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_801 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_800 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_799 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_798 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_797 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_796 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_795 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_794 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_793 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_792 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_791 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_790 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_789 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_788 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_787 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_786 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_785 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_784 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_783 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_782 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_781 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_780 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_779 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_778 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_777 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_776 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_775 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_774 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_773 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_772 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_771 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_770 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_769 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_768 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_767 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_766 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_765 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_764 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_763 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_762 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_761 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_760 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_759 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_758 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_757 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_756 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_755 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_754 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_753 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_752 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_751 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_750 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_749 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_748 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_747 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_746 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_745 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_744 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_743 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_742 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_741 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_740 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_739 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_738 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_737 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_736 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_735 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_734 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_733 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_732 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_731 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_730 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_729 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_728 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_727 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_726 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_725 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_724 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_723 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_722 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_721 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_720 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_719 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_718 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_717 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_716 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_715 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_714 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_713 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_712 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_711 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_710 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_709 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_708 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_707 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_706 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_705 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_704 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_703 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_702 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_701 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_700 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_699 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_698 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_697 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_696 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_695 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_694 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_693 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_692 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_691 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_690 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_689 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_688 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_687 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_686 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_685 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_684 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_683 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_682 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_681 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_680 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_679 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_678 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_677 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_676 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_675 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_674 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_673 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_672 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_671 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_670 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_669 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_668 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_667 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_666 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_665 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_664 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_663 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_662 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_661 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_660 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_659 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_658 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_657 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_656 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_655 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_654 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_653 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_652 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_651 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_650 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_649 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_648 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_647 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_646 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_645 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_644 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_643 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_642 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_641 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_640 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_639 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_638 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_637 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_636 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_635 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_634 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_633 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_632 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_631 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_630 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_629 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_628 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_627 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_626 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_625 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_624 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_623 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_622 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_621 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_620 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_619 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_618 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_617 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_616 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_615 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_614 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_613 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_612 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_611 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_610 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_609 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_608 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_607 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_606 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_605 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_604 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_603 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_602 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_601 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_600 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_599 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_598 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_597 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_596 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_595 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_594 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_593 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_592 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_591 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_590 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_589 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_588 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_587 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_586 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_585 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_584 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_583 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_582 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_581 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_580 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_579 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_578 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_577 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_576 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_575 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_574 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_573 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_572 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_571 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_570 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_569 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_568 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_567 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_566 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_565 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_564 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_563 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_562 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_561 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_560 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_559 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_558 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_557 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_556 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_555 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_554 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_553 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_552 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_551 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_550 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_549 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_548 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_547 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_546 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_545 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_544 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_543 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_542 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_541 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_540 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_539 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_538 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_537 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_536 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_535 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_534 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_533 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_532 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_531 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_530 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_529 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_528 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_527 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_526 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_525 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_524 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_523 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_522 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_521 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_520 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_519 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_518 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_517 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_516 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_515 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_514 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_513 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_512 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_511 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_510 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_509 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_508 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_507 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_506 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_505 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_504 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_503 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_502 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_501 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_500 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_499 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_498 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_497 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_496 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_495 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_494 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_493 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_492 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_491 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_490 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_489 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_488 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_487 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_486 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_485 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_484 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_483 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_482 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_481 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_480 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_479 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_478 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_477 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_476 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_475 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_474 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_473 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_472 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_471 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_470 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_469 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_468 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_467 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_466 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_465 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_464 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_463 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_462 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_461 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_460 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_459 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_458 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_457 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_456 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_455 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_454 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_453 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_452 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_451 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_450 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_449 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_448 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_447 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_446 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_445 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_444 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_443 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_442 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_441 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_440 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_439 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_438 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_437 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_436 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_435 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_434 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_433 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_432 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_431 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_430 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_429 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_428 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_427 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_426 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_425 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_424 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_423 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_422 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_421 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_420 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_419 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_418 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_417 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_416 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_415 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_414 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_413 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_412 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_411 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_410 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_409 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_408 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_407 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_406 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_405 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_404 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_403 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_402 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_401 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_400 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_399 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_398 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_397 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_396 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_395 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_394 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_393 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_392 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_391 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_390 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_389 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_388 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_387 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_386 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_385 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_384 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_383 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_382 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_381 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_380 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_379 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_378 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_377 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_376 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_375 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_374 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_373 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_372 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_371 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_370 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_369 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_368 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_367 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_366 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_365 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_364 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_363 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_362 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_361 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_360 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_359 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_358 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_357 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_356 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_355 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_354 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_353 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_352 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_351 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_350 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_349 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_348 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_347 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_346 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_345 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_344 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_343 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_342 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_341 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_340 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_339 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_338 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_337 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_336 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_335 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_334 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_333 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_332 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_331 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_330 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_329 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_328 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_327 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_326 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_325 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_324 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_323 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_322 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_321 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_320 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_319 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_318 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_317 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_316 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_315 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_314 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_313 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_312 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_311 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_310 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_309 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_308 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_307 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_306 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_305 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_304 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_303 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_302 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_301 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_300 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_299 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_298 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_297 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_296 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_295 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_294 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_293 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_292 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_291 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_290 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_289 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_288 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_287 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_286 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_285 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_284 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_283 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_282 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_281 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_280 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_279 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_278 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_277 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_276 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_275 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_274 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_273 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_272 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_271 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_270 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_269 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_268 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_267 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_266 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_265 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_264 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_263 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_262 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_261 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_260 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_259 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_258 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_257 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_256 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_255 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_254 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_253 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_252 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_251 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_250 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_249 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_248 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_247 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_246 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_245 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_244 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_243 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_242 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_241 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_240 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_239 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_238 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_237 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_236 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_235 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_234 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_233 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_232 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_231 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_230 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_229 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_228 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_227 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_226 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_225 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_224 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_223 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_222 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_221 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_220 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_219 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_218 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_217 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_216 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_215 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_214 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_213 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_212 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_211 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_210 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_209 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_208 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_207 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_206 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_205 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_204 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_203 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_202 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_201 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_200 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_199 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_198 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_197 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_196 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_195 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_194 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_193 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_192 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_191 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_190 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_189 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_188 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_187 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_186 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_185 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_184 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_183 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_182 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_181 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_180 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_179 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_178 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_177 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_176 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_175 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_174 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_173 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_172 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_171 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_170 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_169 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_168 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_167 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_166 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_165 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_164 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_163 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_162 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_161 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_160 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_159 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_158 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_157 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_156 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_155 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_154 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_153 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_152 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_151 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_150 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_149 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_148 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_147 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_146 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_145 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_144 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_143 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_142 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_141 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_140 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_139 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_138 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_137 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_136 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_135 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_134 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_133 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_132 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_131 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_130 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_129 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_128 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_127 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_126 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_125 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_124 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_123 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_122 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_121 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_120 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_119 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_118 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_117 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_116 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_115 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_114 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_113 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_112 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_111 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_110 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_109 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_108 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_107 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_106 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_105 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_104 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_103 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_102 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_101 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_100 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_99 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_98 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_97 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_96 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_95 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_94 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_93 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_92 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_91 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_90 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_89 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_88 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_87 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_86 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_85 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_84 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_83 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_82 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_81 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_80 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_79 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_78 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_77 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_76 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_75 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_74 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_73 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_72 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_71 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_70 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_69 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_68 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_67 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_66 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_65 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_64 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_63 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_62 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_61 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_60 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_59 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_58 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_57 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_56 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_55 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_54 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_53 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_52 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_51 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_50 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_49 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_48 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_47 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_46 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_45 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_44 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_43 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_42 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_41 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_40 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_39 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_38 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_37 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_36 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_35 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_34 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_33 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_32 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_31 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_30 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_29 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_28 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_27 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_26 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_25 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_24 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_23 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_22 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_21 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_20 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_19 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_18 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_17 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_16 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_15 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_14 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_13 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_12 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_11 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_10 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_9 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_8 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_7 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_6 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_5 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_4 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_3 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_2 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X2_1 VDD VSS FILLCELL_X2 
Xxofiller_FILLCELL_X4_2628 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2627 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2626 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2625 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2624 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2623 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2622 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2621 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2620 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2619 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2618 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2617 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2616 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2615 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2614 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2613 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2612 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2611 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2610 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2609 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2608 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2607 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2606 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2605 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2604 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2603 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2602 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2601 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2600 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2599 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2598 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2597 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2596 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2595 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2594 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2593 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2592 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2591 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2590 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2589 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2588 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2587 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2586 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2585 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2584 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2583 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2582 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2581 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2580 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2579 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2578 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2577 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2576 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2575 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2574 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2573 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2572 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2571 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2570 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2569 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2568 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2567 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2566 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2565 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2564 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2563 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2562 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2561 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2560 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2559 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2558 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2557 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2556 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2555 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2554 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2553 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2552 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2551 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2550 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2549 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2548 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2547 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2546 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2545 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2544 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2543 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2542 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2541 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2540 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2539 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2538 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2537 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2536 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2535 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2534 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2533 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2532 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2531 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2530 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2529 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2528 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2527 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2526 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2525 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2524 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2523 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2522 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2521 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2520 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2519 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2518 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2517 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2516 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2515 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2514 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2513 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2512 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2511 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2510 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2509 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2508 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2507 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2506 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2505 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2504 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2503 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2502 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2501 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2500 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2499 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2498 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2497 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2496 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2495 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2494 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2493 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2492 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2491 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2490 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2489 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2488 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2487 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2486 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2485 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2484 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2483 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2482 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2481 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2480 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2479 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2478 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2477 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2476 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2475 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2474 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2473 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2472 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2471 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2470 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2469 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2468 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2467 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2466 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2465 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2464 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2463 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2462 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2461 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2460 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2459 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2458 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2457 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2456 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2455 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2454 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2453 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2452 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2451 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2450 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2449 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2448 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2447 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2446 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2445 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2444 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2443 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2442 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2441 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2440 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2439 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2438 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2437 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2436 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2435 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2434 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2433 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2432 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2431 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2430 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2429 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2428 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2427 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2426 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2425 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2424 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2423 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2422 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2421 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2420 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2419 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2418 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2417 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2416 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2415 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2414 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2413 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2412 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2411 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2410 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2409 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2408 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2407 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2406 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2405 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2404 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2403 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2402 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2401 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2400 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2399 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2398 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2397 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2396 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2395 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2394 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2393 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2392 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2391 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2390 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2389 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2388 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2387 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2386 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2385 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2384 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2383 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2382 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2381 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2380 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2379 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2378 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2377 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2376 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2375 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2374 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2373 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2372 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2371 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2370 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2369 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2368 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2367 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2366 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2365 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2364 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2363 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2362 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2361 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2360 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2359 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2358 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2357 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2356 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2355 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2354 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2353 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2352 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2351 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2350 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2349 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2348 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2347 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2346 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2345 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2344 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2343 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2342 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2341 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2340 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2339 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2338 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2337 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2336 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2335 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2334 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2333 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2332 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2331 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2330 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2329 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2328 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2327 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2326 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2325 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2324 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2323 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2322 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2321 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2320 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2319 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2318 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2317 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2316 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2315 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2314 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2313 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2312 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2311 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2310 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2309 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2308 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2307 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2306 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2305 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2304 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2303 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2302 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2301 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2300 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2299 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2298 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2297 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2296 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2295 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2294 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2293 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2292 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2291 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2290 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2289 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2288 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2287 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2286 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2285 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2284 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2283 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2282 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2281 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2280 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2279 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2278 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2277 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2276 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2275 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2274 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2273 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2272 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2271 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2270 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2269 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2268 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2267 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2266 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2265 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2264 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2263 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2262 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2261 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2260 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2259 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2258 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2257 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2256 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2255 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2254 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2253 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2252 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2251 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2250 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2249 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2248 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2247 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2246 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2245 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2244 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2243 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2242 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2241 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2240 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2239 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2238 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2237 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2236 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2235 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2234 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2233 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2232 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2231 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2230 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2229 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2228 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2227 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2226 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2225 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2224 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2223 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2222 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2221 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2220 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2219 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2218 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2217 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2216 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2215 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2214 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2213 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2212 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2211 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2210 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2209 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2208 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2207 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2206 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2205 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2204 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2203 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2202 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2201 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2200 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2199 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2198 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2197 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2196 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2195 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2194 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2193 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2192 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2191 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2190 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2189 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2188 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2187 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2186 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2185 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2184 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2183 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2182 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2181 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2180 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2179 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2178 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2177 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2176 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2175 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2174 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2173 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2172 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2171 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2170 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2169 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2168 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2167 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2166 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2165 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2164 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2163 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2162 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2161 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2160 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2159 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2158 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2157 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2156 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2155 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2154 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2153 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2152 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2151 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2150 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2149 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2148 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2147 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2146 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2145 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2144 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2143 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2142 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2141 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2140 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2139 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2138 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2137 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2136 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2135 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2134 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2133 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2132 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2131 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2130 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2129 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2128 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2127 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2126 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2125 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2124 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2123 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2122 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2121 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2120 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2119 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2118 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2117 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2116 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2115 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2114 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2113 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2112 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2111 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2110 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2109 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2108 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2107 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2106 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2105 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2104 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2103 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2102 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2101 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2100 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2099 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2098 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2097 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2096 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2095 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2094 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2093 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2092 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2091 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2090 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2089 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2088 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2087 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2086 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2085 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2084 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2083 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2082 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2081 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2080 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2079 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2078 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2077 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2076 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2075 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2074 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2073 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2072 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2071 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2070 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2069 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2068 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2067 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2066 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2065 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2064 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2063 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2062 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2061 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2060 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2059 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2058 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2057 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2056 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2055 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2054 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2053 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2052 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2051 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2050 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2049 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2048 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2047 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2046 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2045 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2044 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2043 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2042 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2041 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2040 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2039 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2038 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2037 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2036 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2035 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2034 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2033 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2032 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2031 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2030 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2029 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2028 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2027 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2026 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2025 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2024 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2023 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2022 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2021 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2020 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2019 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2018 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2017 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2016 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2015 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2014 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2013 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2012 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2011 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2010 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2009 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2008 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2007 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2006 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2005 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2004 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2003 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2002 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2001 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2000 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1999 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1998 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1997 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1996 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1995 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1994 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1993 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1992 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1991 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1990 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1989 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1988 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1987 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1986 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1985 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1984 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1983 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1982 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1981 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1980 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1979 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1978 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1977 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1976 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1975 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1974 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1973 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1972 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1971 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1970 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1969 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1968 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1967 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1966 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1965 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1964 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1963 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1962 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1961 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1960 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1959 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1958 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1957 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1956 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1955 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1954 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1953 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1952 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1951 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1950 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1949 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1948 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1947 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1946 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1945 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1944 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1943 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1942 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1941 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1940 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1939 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1938 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1937 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1936 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1935 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1934 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1933 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1932 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1931 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1930 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1929 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1928 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1927 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1926 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1925 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1924 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1923 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1922 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1921 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1920 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1919 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1918 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1917 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1916 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1915 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1914 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1913 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1912 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1911 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1910 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1909 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1908 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1907 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1906 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1905 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1904 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1903 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1902 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1901 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1900 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1899 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1898 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1897 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1896 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1895 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1894 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1893 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1892 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1891 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1890 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1889 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1888 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1887 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1886 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1885 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1884 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1883 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1882 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1881 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1880 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1879 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1878 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1877 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1876 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1875 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1874 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1873 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1872 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1871 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1870 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1869 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1868 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1867 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1866 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1865 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1864 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1863 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1862 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1861 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1860 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1859 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1858 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1857 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1856 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1855 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1854 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1853 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1852 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1851 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1850 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1849 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1848 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1847 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1846 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1845 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1844 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1843 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1842 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1841 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1840 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1839 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1838 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1837 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1836 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1835 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1834 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1833 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1832 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1831 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1830 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1829 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1828 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1827 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1826 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1825 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1824 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1823 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1822 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1821 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1820 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1819 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1818 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1817 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1816 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1815 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1814 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1813 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1812 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1811 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1810 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1809 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1808 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1807 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1806 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1805 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1804 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1803 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1802 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1801 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1800 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1799 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1798 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1797 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1796 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1795 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1794 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1793 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1792 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1791 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1790 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1789 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1788 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1787 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1786 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1785 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1784 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1783 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1782 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1781 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1780 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1779 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1778 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1777 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1776 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1775 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1774 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1773 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1772 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1771 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1770 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1769 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1768 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1767 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1766 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1765 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1764 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1763 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1762 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1761 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1760 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1759 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1758 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1757 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1756 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1755 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1754 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1753 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1752 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1751 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1750 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1749 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1748 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1747 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1746 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1745 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1744 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1743 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1742 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1741 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1740 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1739 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1738 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1737 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1736 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1735 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1734 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1733 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1732 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1731 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1730 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1729 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1728 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1727 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1726 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1725 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1724 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1723 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1722 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1721 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1720 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1719 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1718 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1717 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1716 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1715 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1714 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1713 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1712 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1711 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1710 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1709 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1708 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1707 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1706 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1705 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1704 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1703 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1702 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1701 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1700 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1699 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1698 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1697 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1696 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1695 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1694 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1693 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1692 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1691 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1690 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1689 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1688 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1687 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1686 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1685 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1684 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1683 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1682 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1681 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1680 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1679 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1678 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1677 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1676 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1675 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1674 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1673 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1672 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1671 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1670 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1669 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1668 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1667 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1666 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1665 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1664 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1663 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1662 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1661 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1660 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1659 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1658 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1657 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1656 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1655 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1654 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1653 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1652 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1651 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1650 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1649 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1648 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1647 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1646 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1645 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1644 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1643 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1642 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1641 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1640 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1639 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1638 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1637 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1636 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1635 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1634 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1633 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1632 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1631 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1630 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1629 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1628 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1627 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1626 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1625 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1624 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1623 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1622 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1621 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1620 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1619 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1618 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1617 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1616 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1615 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1614 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1613 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1612 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1611 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1610 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1609 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1608 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1607 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1606 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1605 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1604 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1603 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1602 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1601 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1600 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1599 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1598 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1597 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1596 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1595 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1594 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1593 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1592 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1591 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1590 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1589 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1588 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1587 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1586 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1585 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1584 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1583 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1582 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1581 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1580 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1579 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1578 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1577 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1576 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1575 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1574 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1573 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1572 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1571 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1570 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1569 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1568 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1567 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1566 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1565 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1564 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1563 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1562 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1561 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1560 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1559 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1558 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1557 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1556 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1555 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1554 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1553 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1552 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1551 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1550 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1549 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1548 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1547 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1546 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1545 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1544 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1543 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1542 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1541 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1540 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1539 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1538 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1537 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1536 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1535 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1534 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1533 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1532 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1531 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1530 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1529 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1528 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1527 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1526 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1525 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1524 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1523 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1522 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1521 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1520 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1519 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1518 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1517 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1516 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1515 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1514 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1513 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1512 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1511 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1510 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1509 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1508 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1507 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1506 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1505 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1504 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1503 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1502 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1501 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1500 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1499 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1498 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1497 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1496 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1495 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1494 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1493 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1492 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1491 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1490 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1489 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1488 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1487 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1486 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1485 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1484 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1483 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1482 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1481 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1480 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1479 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1478 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1477 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1476 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1475 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1474 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1473 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1472 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1471 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1470 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1469 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1468 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1467 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1466 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1465 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1464 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1463 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1462 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1461 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1460 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1459 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1458 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1457 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1456 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1455 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1454 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1453 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1452 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1451 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1450 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1449 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1448 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1447 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1446 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1445 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1444 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1443 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1442 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1441 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1440 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1439 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1438 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1437 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1436 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1435 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1434 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1433 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1432 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1431 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1430 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1429 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1428 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1427 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1426 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1425 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1424 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1423 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1422 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1421 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1420 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1419 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1418 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1417 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1416 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1415 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1414 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1413 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1412 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1411 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1410 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1409 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1408 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1407 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1406 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1405 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1404 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1403 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1402 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1401 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1400 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1399 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1398 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1397 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1396 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1395 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1394 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1393 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1392 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1391 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1390 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1389 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1388 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1387 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1386 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1385 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1384 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1383 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1382 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1381 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1380 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1379 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1378 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1377 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1376 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1375 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1374 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1373 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1372 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1371 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1370 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1369 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1368 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1367 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1366 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1365 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1364 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1363 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1362 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1361 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1360 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1359 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1358 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1357 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1356 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1355 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1354 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1353 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1352 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1351 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1350 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1349 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1348 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1347 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1346 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1345 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1344 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1343 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1342 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1341 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1340 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1339 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1338 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1337 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1336 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1335 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1334 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1333 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1332 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1331 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1330 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1329 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1328 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1327 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1326 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1325 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1324 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1323 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1322 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1321 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1320 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1319 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1318 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1317 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1316 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1315 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1314 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1313 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1312 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1311 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1310 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1309 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1308 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1307 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1306 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1305 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1304 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1303 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1302 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1301 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1300 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1299 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1298 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1297 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1296 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1295 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1294 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1293 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1292 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1291 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1290 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1289 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1288 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1287 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1286 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1285 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1284 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1283 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1282 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1281 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1280 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1279 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1278 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1277 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1276 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1275 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1274 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1273 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1272 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1271 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1270 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1269 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1268 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1267 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1266 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1265 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1264 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1263 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1262 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1261 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1260 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1259 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1258 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1257 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1256 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1255 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1254 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1253 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1252 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1251 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1250 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1249 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1248 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1247 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1246 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1245 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1244 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1243 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1242 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1241 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1240 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1239 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1238 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1237 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1236 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1235 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1234 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1233 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1232 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1231 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1230 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1229 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1228 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1227 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1226 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1225 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1224 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1223 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1222 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1221 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1220 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1219 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1218 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1217 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1216 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1215 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1214 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1213 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1212 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1211 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1210 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1209 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1208 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1207 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1206 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1205 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1204 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1203 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1202 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1201 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1200 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1199 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1198 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1197 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1196 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1195 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1194 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1193 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1192 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1191 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1190 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1189 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1188 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1187 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1186 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1185 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1184 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1183 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1182 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1181 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1180 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1179 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1178 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1177 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1176 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1175 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1174 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1173 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1172 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1171 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1170 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1169 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1168 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1167 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1166 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1165 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1164 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1163 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1162 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1161 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1160 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1159 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1158 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1157 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1156 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1155 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1154 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1153 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1152 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1151 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1150 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1149 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1148 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1147 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1146 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1145 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1144 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1143 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1142 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1141 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1140 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1139 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1138 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1137 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1136 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1135 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1134 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1133 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1132 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1131 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1130 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1129 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1128 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1127 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1126 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1125 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1124 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1123 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1122 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1121 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1120 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1119 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1118 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1117 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1116 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1115 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1114 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1113 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1112 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1111 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1110 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1109 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1108 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1107 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1106 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1105 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1104 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1103 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1102 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1101 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1100 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1099 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1098 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1097 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1096 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1095 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1094 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1093 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1092 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1091 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1090 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1089 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1088 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1087 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1086 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1085 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1084 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1083 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1082 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1081 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1080 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1079 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1078 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1077 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1076 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1075 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1074 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1073 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1072 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1071 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1070 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1069 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1068 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1067 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1066 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1065 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1064 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1063 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1062 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1061 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1060 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1059 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1058 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1057 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1056 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1055 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1054 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1053 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1052 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1051 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1050 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1049 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1048 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1047 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1046 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1045 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1044 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1043 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1042 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1041 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1040 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1039 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1038 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1037 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1036 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1035 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1034 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1033 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1032 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1031 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1030 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1029 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1028 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1027 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1026 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1025 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1024 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1023 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1022 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1021 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1020 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1019 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1018 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1017 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1016 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1015 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1014 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1013 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1012 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1011 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1010 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1009 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1008 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1007 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1006 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1005 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1004 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1003 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1002 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1001 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1000 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_999 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_998 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_997 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_996 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_995 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_994 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_993 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_992 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_991 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_990 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_989 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_988 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_987 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_986 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_985 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_984 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_983 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_982 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_981 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_980 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_979 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_978 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_977 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_976 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_975 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_974 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_973 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_972 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_971 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_970 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_969 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_968 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_967 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_966 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_965 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_964 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_963 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_962 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_961 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_960 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_959 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_958 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_957 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_956 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_955 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_954 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_953 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_952 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_951 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_950 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_949 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_948 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_947 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_946 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_945 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_944 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_943 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_942 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_941 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_940 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_939 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_938 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_937 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_936 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_935 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_934 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_933 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_932 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_931 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_930 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_929 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_928 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_927 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_926 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_925 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_924 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_923 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_922 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_921 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_920 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_919 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_918 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_917 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_916 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_915 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_914 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_913 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_912 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_911 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_910 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_909 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_908 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_907 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_906 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_905 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_904 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_903 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_902 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_901 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_900 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_899 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_898 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_897 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_896 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_895 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_894 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_893 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_892 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_891 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_890 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_889 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_888 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_887 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_886 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_885 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_884 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_883 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_882 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_881 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_880 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_879 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_878 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_877 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_876 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_875 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_874 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_873 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_872 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_871 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_870 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_869 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_868 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_867 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_866 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_865 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_864 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_863 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_862 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_861 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_860 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_859 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_858 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_857 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_856 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_855 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_854 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_853 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_852 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_851 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_850 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_849 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_848 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_847 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_846 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_845 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_844 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_843 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_842 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_841 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_840 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_839 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_838 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_837 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_836 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_835 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_834 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_833 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_832 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_831 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_830 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_829 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_828 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_827 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_826 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_825 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_824 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_823 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_822 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_821 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_820 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_819 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_818 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_817 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_816 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_815 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_814 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_813 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_812 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_811 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_810 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_809 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_808 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_807 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_806 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_805 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_804 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_803 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_802 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_801 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_800 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_799 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_798 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_797 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_796 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_795 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_794 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_793 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_792 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_791 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_790 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_789 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_788 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_787 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_786 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_785 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_784 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_783 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_782 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_781 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_780 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_779 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_778 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_777 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_776 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_775 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_774 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_773 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_772 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_771 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_770 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_769 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_768 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_767 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_766 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_765 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_764 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_763 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_762 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_761 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_760 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_759 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_758 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_757 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_756 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_755 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_754 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_753 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_752 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_751 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_750 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_749 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_748 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_747 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_746 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_745 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_744 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_743 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_742 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_741 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_740 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_739 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_738 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_737 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_736 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_735 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_734 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_733 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_732 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_731 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_730 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_729 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_728 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_727 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_726 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_725 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_724 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_723 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_722 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_721 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_720 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_719 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_718 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_717 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_716 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_715 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_714 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_713 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_712 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_711 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_710 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_709 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_708 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_707 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_706 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_705 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_704 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_703 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_702 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_701 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_700 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_699 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_698 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_697 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_696 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_695 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_694 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_693 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_692 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_691 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_690 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_689 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_688 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_687 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_686 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_685 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_684 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_683 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_682 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_681 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_680 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_679 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_678 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_677 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_676 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_675 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_674 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_673 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_672 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_671 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_670 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_669 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_668 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_667 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_666 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_665 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_664 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_663 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_662 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_661 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_660 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_659 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_658 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_657 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_656 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_655 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_654 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_653 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_652 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_651 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_650 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_649 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_648 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_647 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_646 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_645 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_644 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_643 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_642 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_641 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_640 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_639 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_638 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_637 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_636 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_635 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_634 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_633 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_632 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_631 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_630 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_629 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_628 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_627 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_626 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_625 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_624 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_623 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_622 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_621 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_620 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_619 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_618 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_617 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_616 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_615 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_614 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_613 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_612 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_611 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_610 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_609 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_608 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_607 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_606 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_605 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_604 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_603 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_602 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_601 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_600 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_599 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_598 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_597 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_596 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_595 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_594 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_593 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_592 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_591 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_590 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_589 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_588 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_587 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_586 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_585 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_584 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_583 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_582 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_581 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_580 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_579 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_578 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_577 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_576 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_575 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_574 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_573 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_572 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_571 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_570 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_569 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_568 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_567 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_566 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_565 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_564 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_563 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_562 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_561 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_560 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_559 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_558 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_557 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_556 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_555 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_554 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_553 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_552 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_551 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_550 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_549 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_548 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_547 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_546 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_545 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_544 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_543 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_542 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_541 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_540 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_539 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_538 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_537 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_536 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_535 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_534 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_533 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_532 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_531 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_530 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_529 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_528 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_527 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_526 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_525 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_524 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_523 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_522 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_521 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_520 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_519 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_518 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_517 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_516 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_515 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_514 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_513 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_512 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_511 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_510 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_509 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_508 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_507 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_506 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_505 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_504 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_503 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_502 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_501 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_500 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_499 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_498 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_497 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_496 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_495 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_494 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_493 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_492 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_491 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_490 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_489 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_488 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_487 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_486 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_485 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_484 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_483 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_482 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_481 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_480 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_479 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_478 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_477 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_476 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_475 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_474 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_473 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_472 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_471 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_470 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_469 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_468 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_467 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_466 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_465 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_464 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_463 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_462 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_461 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_460 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_459 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_458 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_457 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_456 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_455 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_454 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_453 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_452 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_451 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_450 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_449 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_448 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_447 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_446 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_445 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_444 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_443 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_442 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_441 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_440 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_439 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_438 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_437 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_436 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_435 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_434 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_433 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_432 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_431 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_430 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_429 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_428 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_427 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_426 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_425 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_424 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_423 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_422 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_421 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_420 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_419 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_418 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_417 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_416 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_415 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_414 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_413 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_412 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_411 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_410 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_409 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_408 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_407 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_406 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_405 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_404 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_403 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_402 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_401 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_400 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_399 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_398 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_397 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_396 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_395 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_394 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_393 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_392 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_391 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_390 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_389 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_388 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_387 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_386 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_385 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_384 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_383 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_382 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_381 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_380 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_379 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_378 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_377 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_376 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_375 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_374 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_373 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_372 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_371 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_370 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_369 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_368 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_367 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_366 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_365 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_364 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_363 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_362 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_361 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_360 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_359 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_358 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_357 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_356 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_355 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_354 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_353 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_352 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_351 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_350 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_349 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_348 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_347 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_346 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_345 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_344 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_343 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_342 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_341 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_340 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_339 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_338 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_337 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_336 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_335 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_334 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_333 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_332 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_331 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_330 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_329 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_328 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_327 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_326 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_325 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_324 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_323 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_322 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_321 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_320 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_319 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_318 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_317 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_316 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_315 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_314 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_313 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_312 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_311 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_310 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_309 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_308 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_307 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_306 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_305 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_304 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_303 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_302 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_301 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_300 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_299 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_298 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_297 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_296 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_295 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_294 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_293 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_292 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_291 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_290 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_289 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_288 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_287 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_286 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_285 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_284 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_283 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_282 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_281 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_280 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_279 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_278 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_277 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_276 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_275 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_274 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_273 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_272 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_271 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_270 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_269 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_268 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_267 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_266 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_265 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_264 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_263 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_262 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_261 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_260 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_259 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_258 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_257 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_256 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_255 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_254 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_253 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_252 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_251 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_250 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_249 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_248 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_247 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_246 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_245 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_244 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_243 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_242 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_241 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_240 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_239 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_238 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_237 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_236 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_235 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_234 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_233 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_232 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_231 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_230 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_229 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_228 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_227 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_226 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_225 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_224 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_223 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_222 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_221 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_220 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_219 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_218 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_217 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_216 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_215 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_214 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_213 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_212 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_211 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_210 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_209 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_208 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_207 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_206 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_205 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_204 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_203 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_202 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_201 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_200 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_199 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_198 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_197 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_196 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_195 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_194 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_193 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_192 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_191 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_190 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_189 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_188 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_187 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_186 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_185 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_184 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_183 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_182 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_181 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_180 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_179 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_178 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_177 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_176 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_175 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_174 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_173 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_172 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_171 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_170 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_169 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_168 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_167 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_166 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_165 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_164 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_163 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_162 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_161 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_160 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_159 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_158 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_157 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_156 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_155 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_154 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_153 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_152 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_151 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_150 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_149 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_148 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_147 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_146 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_145 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_144 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_143 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_142 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_141 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_140 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_139 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_138 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_137 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_136 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_135 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_134 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_133 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_132 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_131 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_130 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_129 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_128 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_127 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_126 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_125 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_124 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_123 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_122 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_121 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_120 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_119 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_118 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_117 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_116 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_115 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_114 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_113 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_112 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_111 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_110 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_109 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_108 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_107 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_106 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_105 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_104 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_103 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_102 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_101 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_100 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_99 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_98 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_97 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_96 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_95 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_94 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_93 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_92 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_91 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_90 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_89 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_88 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_87 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_86 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_85 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_84 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_83 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_82 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_81 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_80 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_79 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_78 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_77 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_76 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_75 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_74 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_73 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_72 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_71 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_70 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_69 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_68 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_67 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_66 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_65 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_64 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_63 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_62 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_61 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_60 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_59 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_58 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_57 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_56 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_55 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_54 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_53 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_52 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_51 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_50 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_49 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_48 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_47 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_46 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_45 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_44 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_43 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_42 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_41 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_40 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_39 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_38 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_37 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_36 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_35 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_34 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_33 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_32 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_31 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_30 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_29 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_28 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_27 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_26 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_25 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_24 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_23 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_22 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_21 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_20 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_19 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_18 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_17 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_16 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_15 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_14 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_13 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_12 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_11 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_10 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_9 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_8 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_7 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_6 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_5 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_4 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_3 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_2 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X4_1 VDD VSS FILLCELL_X4 
Xxofiller_FILLCELL_X8_2260 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2259 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2258 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2257 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2256 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2255 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2254 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2253 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2252 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2251 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2250 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2249 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2248 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2247 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2246 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2245 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2244 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2243 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2242 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2241 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2240 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2239 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2238 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2237 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2236 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2235 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2234 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2233 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2232 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2231 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2230 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2229 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2228 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2227 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2226 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2225 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2224 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2223 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2222 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2221 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2220 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2219 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2218 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2217 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2216 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2215 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2214 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2213 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2212 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2211 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2210 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2209 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2208 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2207 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2206 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2205 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2204 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2203 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2202 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2201 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2200 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2199 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2198 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2197 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2196 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2195 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2194 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2193 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2192 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2191 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2190 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2189 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2188 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2187 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2186 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2185 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2184 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2183 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2182 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2181 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2180 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2179 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2178 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2177 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2176 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2175 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2174 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2173 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2172 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2171 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2170 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2169 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2168 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2167 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2166 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2165 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2164 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2163 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2162 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2161 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2160 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2159 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2158 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2157 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2156 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2155 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2154 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2153 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2152 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2151 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2150 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2149 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2148 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2147 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2146 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2145 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2144 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2143 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2142 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2141 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2140 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2139 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2138 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2137 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2136 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2135 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2134 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2133 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2132 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2131 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2130 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2129 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2128 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2127 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2126 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2125 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2124 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2123 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2122 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2121 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2120 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2119 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2118 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2117 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2116 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2115 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2114 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2113 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2112 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2111 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2110 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2109 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2108 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2107 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2106 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2105 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2104 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2103 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2102 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2101 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2100 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2099 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2098 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2097 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2096 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2095 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2094 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2093 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2092 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2091 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2090 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2089 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2088 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2087 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2086 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2085 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2084 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2083 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2082 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2081 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2080 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2079 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2078 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2077 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2076 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2075 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2074 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2073 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2072 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2071 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2070 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2069 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2068 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2067 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2066 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2065 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2064 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2063 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2062 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2061 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2060 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2059 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2058 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2057 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2056 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2055 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2054 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2053 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2052 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2051 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2050 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2049 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2048 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2047 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2046 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2045 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2044 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2043 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2042 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2041 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2040 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2039 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2038 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2037 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2036 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2035 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2034 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2033 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2032 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2031 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2030 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2029 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2028 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2027 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2026 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2025 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2024 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2023 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2022 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2021 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2020 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2019 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2018 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2017 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2016 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2015 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2014 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2013 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2012 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2011 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2010 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2009 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2008 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2007 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2006 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2005 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2004 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2003 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2002 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2001 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2000 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1999 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1998 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1997 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1996 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1995 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1994 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1993 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1992 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1991 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1990 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1989 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1988 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1987 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1986 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1985 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1984 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1983 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1982 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1981 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1980 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1979 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1978 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1977 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1976 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1975 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1974 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1973 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1972 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1971 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1970 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1969 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1968 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1967 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1966 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1965 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1964 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1963 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1962 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1961 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1960 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1959 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1958 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1957 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1956 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1955 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1954 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1953 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1952 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1951 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1950 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1949 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1948 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1947 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1946 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1945 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1944 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1943 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1942 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1941 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1940 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1939 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1938 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1937 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1936 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1935 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1934 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1933 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1932 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1931 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1930 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1929 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1928 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1927 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1926 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1925 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1924 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1923 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1922 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1921 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1920 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1919 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1918 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1917 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1916 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1915 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1914 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1913 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1912 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1911 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1910 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1909 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1908 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1907 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1906 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1905 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1904 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1903 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1902 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1901 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1900 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1899 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1898 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1897 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1896 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1895 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1894 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1893 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1892 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1891 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1890 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1889 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1888 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1887 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1886 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1885 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1884 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1883 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1882 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1881 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1880 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1879 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1878 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1877 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1876 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1875 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1874 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1873 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1872 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1871 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1870 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1869 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1868 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1867 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1866 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1865 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1864 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1863 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1862 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1861 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1860 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1859 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1858 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1857 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1856 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1855 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1854 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1853 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1852 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1851 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1850 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1849 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1848 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1847 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1846 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1845 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1844 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1843 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1842 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1841 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1840 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1839 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1838 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1837 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1836 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1835 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1834 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1833 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1832 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1831 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1830 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1829 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1828 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1827 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1826 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1825 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1824 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1823 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1822 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1821 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1820 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1819 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1818 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1817 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1816 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1815 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1814 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1813 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1812 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1811 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1810 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1809 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1808 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1807 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1806 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1805 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1804 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1803 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1802 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1801 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1800 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1799 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1798 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1797 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1796 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1795 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1794 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1793 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1792 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1791 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1790 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1789 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1788 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1787 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1786 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1785 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1784 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1783 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1782 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1781 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1780 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1779 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1778 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1777 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1776 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1775 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1774 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1773 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1772 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1771 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1770 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1769 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1768 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1767 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1766 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1765 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1764 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1763 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1762 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1761 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1760 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1759 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1758 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1757 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1756 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1755 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1754 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1753 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1752 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1751 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1750 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1749 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1748 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1747 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1746 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1745 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1744 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1743 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1742 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1741 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1740 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1739 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1738 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1737 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1736 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1735 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1734 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1733 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1732 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1731 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1730 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1729 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1728 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1727 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1726 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1725 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1724 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1723 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1722 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1721 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1720 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1719 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1718 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1717 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1716 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1715 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1714 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1713 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1712 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1711 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1710 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1709 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1708 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1707 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1706 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1705 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1704 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1703 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1702 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1701 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1700 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1699 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1698 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1697 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1696 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1695 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1694 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1693 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1692 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1691 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1690 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1689 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1688 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1687 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1686 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1685 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1684 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1683 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1682 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1681 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1680 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1679 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1678 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1677 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1676 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1675 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1674 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1673 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1672 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1671 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1670 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1669 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1668 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1667 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1666 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1665 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1664 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1663 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1662 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1661 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1660 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1659 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1658 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1657 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1656 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1655 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1654 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1653 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1652 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1651 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1650 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1649 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1648 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1647 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1646 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1645 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1644 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1643 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1642 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1641 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1640 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1639 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1638 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1637 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1636 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1635 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1634 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1633 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1632 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1631 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1630 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1629 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1628 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1627 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1626 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1625 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1624 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1623 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1622 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1621 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1620 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1619 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1618 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1617 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1616 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1615 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1614 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1613 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1612 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1611 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1610 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1609 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1608 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1607 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1606 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1605 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1604 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1603 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1602 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1601 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1600 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1599 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1598 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1597 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1596 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1595 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1594 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1593 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1592 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1591 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1590 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1589 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1588 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1587 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1586 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1585 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1584 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1583 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1582 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1581 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1580 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1579 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1578 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1577 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1576 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1575 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1574 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1573 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1572 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1571 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1570 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1569 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1568 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1567 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1566 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1565 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1564 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1563 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1562 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1561 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1560 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1559 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1558 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1557 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1556 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1555 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1554 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1553 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1552 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1551 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1550 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1549 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1548 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1547 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1546 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1545 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1544 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1543 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1542 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1541 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1540 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1539 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1538 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1537 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1536 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1535 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1534 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1533 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1532 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1531 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1530 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1529 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1528 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1527 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1526 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1525 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1524 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1523 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1522 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1521 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1520 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1519 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1518 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1517 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1516 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1515 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1514 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1513 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1512 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1511 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1510 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1509 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1508 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1507 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1506 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1505 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1504 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1503 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1502 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1501 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1500 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1499 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1498 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1497 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1496 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1495 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1494 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1493 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1492 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1491 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1490 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1489 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1488 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1487 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1486 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1485 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1484 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1483 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1482 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1481 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1480 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1479 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1478 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1477 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1476 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1475 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1474 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1473 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1472 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1471 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1470 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1469 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1468 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1467 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1466 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1465 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1464 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1463 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1462 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1461 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1460 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1459 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1458 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1457 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1456 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1455 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1454 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1453 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1452 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1451 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1450 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1449 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1448 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1447 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1446 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1445 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1444 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1443 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1442 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1441 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1440 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1439 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1438 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1437 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1436 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1435 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1434 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1433 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1432 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1431 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1430 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1429 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1428 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1427 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1426 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1425 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1424 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1423 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1422 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1421 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1420 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1419 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1418 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1417 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1416 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1415 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1414 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1413 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1412 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1411 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1410 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1409 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1408 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1407 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1406 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1405 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1404 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1403 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1402 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1401 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1400 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1399 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1398 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1397 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1396 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1395 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1394 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1393 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1392 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1391 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1390 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1389 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1388 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1387 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1386 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1385 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1384 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1383 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1382 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1381 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1380 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1379 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1378 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1377 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1376 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1375 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1374 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1373 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1372 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1371 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1370 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1369 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1368 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1367 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1366 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1365 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1364 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1363 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1362 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1361 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1360 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1359 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1358 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1357 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1356 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1355 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1354 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1353 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1352 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1351 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1350 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1349 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1348 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1347 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1346 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1345 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1344 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1343 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1342 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1341 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1340 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1339 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1338 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1337 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1336 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1335 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1334 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1333 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1332 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1331 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1330 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1329 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1328 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1327 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1326 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1325 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1324 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1323 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1322 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1321 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1320 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1319 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1318 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1317 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1316 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1315 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1314 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1313 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1312 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1311 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1310 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1309 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1308 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1307 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1306 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1305 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1304 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1303 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1302 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1301 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1300 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1299 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1298 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1297 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1296 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1295 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1294 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1293 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1292 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1291 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1290 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1289 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1288 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1287 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1286 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1285 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1284 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1283 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1282 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1281 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1280 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1279 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1278 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1277 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1276 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1275 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1274 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1273 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1272 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1271 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1270 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1269 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1268 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1267 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1266 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1265 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1264 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1263 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1262 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1261 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1260 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1259 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1258 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1257 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1256 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1255 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1254 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1253 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1252 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1251 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1250 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1249 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1248 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1247 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1246 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1245 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1244 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1243 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1242 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1241 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1240 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1239 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1238 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1237 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1236 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1235 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1234 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1233 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1232 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1231 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1230 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1229 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1228 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1227 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1226 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1225 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1224 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1223 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1222 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1221 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1220 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1219 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1218 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1217 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1216 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1215 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1214 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1213 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1212 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1211 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1210 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1209 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1208 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1207 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1206 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1205 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1204 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1203 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1202 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1201 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1200 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1199 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1198 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1197 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1196 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1195 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1194 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1193 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1192 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1191 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1190 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1189 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1188 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1187 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1186 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1185 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1184 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1183 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1182 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1181 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1180 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1179 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1178 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1177 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1176 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1175 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1174 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1173 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1172 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1171 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1170 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1169 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1168 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1167 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1166 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1165 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1164 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1163 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1162 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1161 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1160 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1159 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1158 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1157 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1156 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1155 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1154 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1153 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1152 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1151 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1150 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1149 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1148 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1147 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1146 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1145 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1144 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1143 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1142 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1141 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1140 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1139 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1138 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1137 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1136 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1135 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1134 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1133 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1132 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1131 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1130 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1129 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1128 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1127 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1126 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1125 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1124 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1123 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1122 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1121 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1120 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1119 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1118 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1117 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1116 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1115 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1114 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1113 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1112 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1111 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1110 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1109 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1108 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1107 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1106 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1105 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1104 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1103 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1102 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1101 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1100 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1099 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1098 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1097 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1096 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1095 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1094 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1093 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1092 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1091 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1090 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1089 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1088 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1087 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1086 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1085 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1084 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1083 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1082 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1081 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1080 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1079 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1078 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1077 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1076 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1075 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1074 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1073 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1072 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1071 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1070 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1069 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1068 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1067 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1066 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1065 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1064 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1063 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1062 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1061 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1060 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1059 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1058 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1057 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1056 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1055 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1054 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1053 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1052 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1051 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1050 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1049 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1048 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1047 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1046 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1045 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1044 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1043 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1042 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1041 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1040 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1039 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1038 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1037 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1036 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1035 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1034 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1033 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1032 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1031 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1030 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1029 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1028 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1027 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1026 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1025 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1024 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1023 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1022 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1021 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1020 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1019 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1018 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1017 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1016 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1015 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1014 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1013 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1012 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1011 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1010 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1009 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1008 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1007 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1006 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1005 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1004 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1003 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1002 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1001 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1000 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_999 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_998 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_997 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_996 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_995 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_994 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_993 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_992 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_991 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_990 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_989 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_988 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_987 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_986 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_985 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_984 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_983 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_982 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_981 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_980 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_979 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_978 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_977 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_976 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_975 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_974 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_973 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_972 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_971 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_970 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_969 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_968 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_967 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_966 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_965 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_964 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_963 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_962 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_961 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_960 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_959 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_958 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_957 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_956 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_955 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_954 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_953 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_952 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_951 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_950 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_949 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_948 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_947 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_946 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_945 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_944 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_943 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_942 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_941 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_940 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_939 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_938 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_937 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_936 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_935 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_934 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_933 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_932 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_931 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_930 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_929 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_928 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_927 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_926 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_925 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_924 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_923 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_922 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_921 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_920 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_919 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_918 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_917 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_916 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_915 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_914 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_913 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_912 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_911 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_910 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_909 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_908 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_907 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_906 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_905 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_904 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_903 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_902 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_901 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_900 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_899 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_898 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_897 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_896 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_895 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_894 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_893 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_892 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_891 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_890 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_889 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_888 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_887 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_886 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_885 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_884 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_883 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_882 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_881 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_880 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_879 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_878 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_877 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_876 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_875 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_874 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_873 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_872 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_871 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_870 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_869 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_868 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_867 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_866 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_865 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_864 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_863 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_862 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_861 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_860 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_859 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_858 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_857 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_856 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_855 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_854 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_853 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_852 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_851 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_850 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_849 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_848 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_847 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_846 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_845 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_844 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_843 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_842 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_841 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_840 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_839 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_838 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_837 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_836 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_835 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_834 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_833 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_832 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_831 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_830 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_829 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_828 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_827 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_826 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_825 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_824 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_823 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_822 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_821 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_820 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_819 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_818 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_817 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_816 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_815 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_814 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_813 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_812 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_811 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_810 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_809 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_808 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_807 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_806 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_805 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_804 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_803 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_802 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_801 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_800 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_799 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_798 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_797 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_796 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_795 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_794 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_793 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_792 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_791 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_790 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_789 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_788 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_787 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_786 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_785 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_784 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_783 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_782 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_781 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_780 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_779 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_778 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_777 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_776 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_775 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_774 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_773 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_772 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_771 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_770 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_769 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_768 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_767 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_766 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_765 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_764 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_763 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_762 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_761 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_760 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_759 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_758 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_757 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_756 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_755 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_754 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_753 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_752 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_751 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_750 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_749 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_748 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_747 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_746 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_745 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_744 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_743 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_742 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_741 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_740 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_739 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_738 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_737 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_736 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_735 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_734 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_733 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_732 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_731 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_730 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_729 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_728 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_727 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_726 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_725 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_724 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_723 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_722 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_721 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_720 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_719 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_718 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_717 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_716 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_715 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_714 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_713 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_712 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_711 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_710 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_709 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_708 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_707 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_706 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_705 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_704 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_703 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_702 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_701 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_700 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_699 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_698 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_697 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_696 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_695 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_694 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_693 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_692 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_691 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_690 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_689 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_688 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_687 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_686 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_685 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_684 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_683 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_682 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_681 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_680 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_679 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_678 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_677 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_676 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_675 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_674 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_673 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_672 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_671 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_670 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_669 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_668 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_667 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_666 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_665 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_664 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_663 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_662 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_661 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_660 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_659 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_658 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_657 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_656 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_655 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_654 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_653 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_652 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_651 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_650 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_649 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_648 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_647 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_646 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_645 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_644 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_643 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_642 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_641 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_640 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_639 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_638 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_637 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_636 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_635 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_634 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_633 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_632 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_631 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_630 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_629 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_628 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_627 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_626 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_625 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_624 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_623 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_622 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_621 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_620 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_619 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_618 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_617 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_616 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_615 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_614 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_613 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_612 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_611 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_610 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_609 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_608 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_607 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_606 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_605 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_604 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_603 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_602 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_601 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_600 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_599 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_598 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_597 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_596 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_595 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_594 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_593 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_592 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_591 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_590 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_589 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_588 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_587 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_586 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_585 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_584 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_583 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_582 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_581 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_580 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_579 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_578 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_577 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_576 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_575 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_574 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_573 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_572 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_571 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_570 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_569 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_568 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_567 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_566 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_565 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_564 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_563 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_562 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_561 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_560 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_559 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_558 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_557 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_556 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_555 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_554 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_553 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_552 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_551 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_550 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_549 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_548 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_547 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_546 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_545 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_544 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_543 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_542 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_541 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_540 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_539 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_538 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_537 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_536 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_535 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_534 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_533 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_532 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_531 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_530 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_529 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_528 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_527 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_526 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_525 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_524 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_523 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_522 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_521 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_520 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_519 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_518 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_517 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_516 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_515 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_514 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_513 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_512 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_511 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_510 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_509 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_508 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_507 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_506 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_505 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_504 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_503 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_502 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_501 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_500 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_499 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_498 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_497 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_496 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_495 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_494 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_493 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_492 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_491 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_490 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_489 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_488 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_487 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_486 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_485 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_484 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_483 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_482 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_481 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_480 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_479 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_478 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_477 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_476 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_475 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_474 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_473 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_472 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_471 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_470 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_469 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_468 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_467 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_466 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_465 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_464 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_463 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_462 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_461 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_460 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_459 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_458 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_457 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_456 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_455 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_454 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_453 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_452 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_451 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_450 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_449 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_448 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_447 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_446 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_445 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_444 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_443 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_442 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_441 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_440 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_439 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_438 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_437 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_436 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_435 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_434 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_433 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_432 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_431 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_430 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_429 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_428 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_427 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_426 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_425 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_424 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_423 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_422 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_421 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_420 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_419 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_418 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_417 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_416 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_415 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_414 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_413 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_412 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_411 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_410 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_409 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_408 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_407 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_406 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_405 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_404 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_403 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_402 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_401 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_400 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_399 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_398 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_397 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_396 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_395 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_394 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_393 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_392 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_391 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_390 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_389 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_388 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_387 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_386 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_385 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_384 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_383 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_382 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_381 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_380 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_379 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_378 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_377 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_376 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_375 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_374 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_373 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_372 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_371 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_370 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_369 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_368 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_367 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_366 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_365 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_364 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_363 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_362 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_361 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_360 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_359 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_358 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_357 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_356 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_355 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_354 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_353 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_352 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_351 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_350 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_349 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_348 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_347 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_346 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_345 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_344 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_343 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_342 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_341 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_340 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_339 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_338 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_337 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_336 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_335 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_334 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_333 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_332 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_331 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_330 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_329 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_328 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_327 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_326 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_325 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_324 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_323 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_322 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_321 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_320 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_319 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_318 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_317 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_316 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_315 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_314 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_313 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_312 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_311 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_310 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_309 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_308 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_307 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_306 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_305 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_304 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_303 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_302 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_301 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_300 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_299 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_298 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_297 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_296 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_295 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_294 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_293 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_292 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_291 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_290 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_289 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_288 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_287 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_286 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_285 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_284 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_283 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_282 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_281 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_280 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_279 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_278 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_277 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_276 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_275 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_274 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_273 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_272 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_271 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_270 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_269 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_268 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_267 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_266 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_265 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_264 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_263 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_262 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_261 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_260 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_259 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_258 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_257 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_256 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_255 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_254 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_253 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_252 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_251 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_250 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_249 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_248 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_247 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_246 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_245 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_244 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_243 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_242 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_241 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_240 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_239 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_238 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_237 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_236 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_235 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_234 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_233 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_232 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_231 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_230 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_229 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_228 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_227 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_226 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_225 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_224 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_223 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_222 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_221 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_220 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_219 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_218 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_217 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_216 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_215 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_214 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_213 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_212 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_211 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_210 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_209 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_208 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_207 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_206 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_205 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_204 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_203 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_202 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_201 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_200 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_199 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_198 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_197 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_196 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_195 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_194 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_193 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_192 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_191 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_190 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_189 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_188 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_187 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_186 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_185 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_184 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_183 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_182 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_181 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_180 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_179 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_178 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_177 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_176 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_175 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_174 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_173 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_172 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_171 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_170 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_169 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_168 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_167 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_166 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_165 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_164 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_163 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_162 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_161 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_160 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_159 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_158 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_157 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_156 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_155 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_154 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_153 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_152 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_151 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_150 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_149 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_148 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_147 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_146 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_145 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_144 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_143 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_142 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_141 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_140 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_139 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_138 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_137 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_136 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_135 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_134 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_133 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_132 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_131 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_130 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_129 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_128 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_127 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_126 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_125 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_124 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_123 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_122 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_121 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_120 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_119 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_118 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_117 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_116 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_115 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_114 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_113 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_112 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_111 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_110 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_109 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_108 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_107 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_106 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_105 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_104 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_103 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_102 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_101 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_100 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_99 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_98 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_97 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_96 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_95 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_94 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_93 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_92 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_91 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_90 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_89 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_88 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_87 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_86 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_85 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_84 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_83 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_82 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_81 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_80 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_79 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_78 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_77 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_76 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_75 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_74 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_73 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_72 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_71 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_70 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_69 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_68 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_67 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_66 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_65 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_64 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_63 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_62 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_61 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_60 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_59 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_58 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_57 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_56 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_55 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_54 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_53 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_52 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_51 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_50 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_49 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_48 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_47 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_46 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_45 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_44 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_43 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_42 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_41 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_40 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_39 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_38 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_37 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_36 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_35 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_34 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_33 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_32 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_31 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_30 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_29 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_28 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_27 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_26 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_25 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_24 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_23 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_22 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_21 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_20 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_19 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_18 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_17 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_16 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_15 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_14 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_13 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_12 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_11 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_10 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_9 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_8 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_7 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_6 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_5 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_4 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_3 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_2 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X8_1 VDD VSS FILLCELL_X8 
Xxofiller_FILLCELL_X16_999 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_998 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_997 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_996 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_995 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_994 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_993 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_992 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_991 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_990 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_989 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_988 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_987 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_986 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_985 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_984 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_983 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_982 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_981 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_980 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_979 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_978 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_977 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_976 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_975 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_974 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_973 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_972 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_971 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_970 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_969 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_968 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_967 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_966 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_965 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_964 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_963 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_962 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_961 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_960 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_959 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_958 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_957 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_956 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_955 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_954 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_953 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_952 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_951 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_950 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_949 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_948 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_947 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_946 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_945 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_944 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_943 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_942 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_941 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_940 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_939 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_938 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_937 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_936 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_935 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_934 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_933 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_932 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_931 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_930 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_929 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_928 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_927 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_926 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_925 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_924 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_923 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_922 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_921 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_920 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_919 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_918 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_917 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_916 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_915 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_914 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_913 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_912 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_911 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_910 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_909 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_908 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_907 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_906 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_905 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_904 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_903 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_902 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_901 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_900 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_899 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_898 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_897 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_896 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_895 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_894 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_893 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_892 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_891 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_890 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_889 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_888 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_887 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_886 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_885 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_884 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_883 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_882 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_881 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_880 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_879 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_878 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_877 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_876 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_875 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_874 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_873 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_872 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_871 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_870 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_869 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_868 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_867 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_866 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_865 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_864 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_863 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_862 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_861 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_860 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_859 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_858 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_857 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_856 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_855 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_854 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_853 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_852 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_851 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_850 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_849 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_848 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_847 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_846 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_845 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_844 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_843 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_842 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_841 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_840 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_839 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_838 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_837 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_836 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_835 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_834 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_833 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_832 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_831 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_830 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_829 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_828 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_827 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_826 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_825 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_824 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_823 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_822 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_821 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_820 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_819 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_818 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_817 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_816 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_815 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_814 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_813 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_812 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_811 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_810 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_809 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_808 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_807 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_806 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_805 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_804 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_803 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_802 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_801 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_800 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_799 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_798 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_797 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_796 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_795 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_794 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_793 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_792 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_791 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_790 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_789 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_788 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_787 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_786 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_785 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_784 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_783 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_782 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_781 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_780 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_779 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_778 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_777 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_776 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_775 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_774 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_773 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_772 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_771 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_770 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_769 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_768 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_767 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_766 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_765 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_764 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_763 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_762 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_761 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_760 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_759 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_758 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_757 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_756 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_755 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_754 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_753 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_752 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_751 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_750 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_749 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_748 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_747 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_746 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_745 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_744 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_743 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_742 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_741 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_740 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_739 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_738 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_737 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_736 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_735 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_734 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_733 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_732 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_731 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_730 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_729 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_728 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_727 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_726 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_725 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_724 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_723 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_722 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_721 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_720 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_719 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_718 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_717 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_716 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_715 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_714 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_713 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_712 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_711 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_710 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_709 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_708 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_707 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_706 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_705 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_704 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_703 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_702 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_701 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_700 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_699 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_698 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_697 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_696 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_695 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_694 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_693 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_692 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_691 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_690 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_689 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_688 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_687 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_686 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_685 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_684 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_683 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_682 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_681 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_680 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_679 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_678 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_677 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_676 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_675 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_674 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_673 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_672 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_671 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_670 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_669 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_668 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_667 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_666 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_665 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_664 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_663 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_662 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_661 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_660 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_659 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_658 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_657 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_656 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_655 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_654 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_653 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_652 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_651 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_650 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_649 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_648 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_647 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_646 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_645 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_644 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_643 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_642 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_641 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_640 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_639 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_638 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_637 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_636 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_635 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_634 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_633 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_632 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_631 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_630 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_629 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_628 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_627 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_626 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_625 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_624 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_623 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_622 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_621 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_620 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_619 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_618 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_617 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_616 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_615 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_614 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_613 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_612 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_611 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_610 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_609 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_608 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_607 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_606 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_605 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_604 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_603 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_602 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_601 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_600 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_599 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_598 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_597 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_596 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_595 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_594 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_593 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_592 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_591 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_590 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_589 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_588 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_587 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_586 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_585 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_584 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_583 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_582 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_581 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_580 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_579 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_578 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_577 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_576 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_575 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_574 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_573 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_572 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_571 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_570 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_569 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_568 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_567 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_566 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_565 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_564 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_563 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_562 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_561 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_560 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_559 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_558 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_557 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_556 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_555 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_554 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_553 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_552 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_551 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_550 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_549 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_548 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_547 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_546 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_545 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_544 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_543 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_542 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_541 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_540 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_539 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_538 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_537 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_536 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_535 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_534 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_533 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_532 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_531 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_530 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_529 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_528 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_527 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_526 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_525 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_524 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_523 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_522 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_521 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_520 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_519 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_518 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_517 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_516 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_515 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_514 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_513 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_512 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_511 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_510 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_509 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_508 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_507 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_506 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_505 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_504 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_503 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_502 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_501 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_500 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_499 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_498 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_497 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_496 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_495 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_494 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_493 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_492 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_491 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_490 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_489 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_488 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_487 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_486 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_485 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_484 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_483 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_482 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_481 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_480 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_479 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_478 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_477 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_476 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_475 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_474 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_473 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_472 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_471 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_470 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_469 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_468 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_467 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_466 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_465 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_464 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_463 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_462 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_461 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_460 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_459 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_458 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_457 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_456 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_455 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_454 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_453 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_452 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_451 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_450 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_449 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_448 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_447 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_446 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_445 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_444 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_443 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_442 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_441 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_440 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_439 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_438 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_437 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_436 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_435 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_434 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_433 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_432 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_431 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_430 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_429 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_428 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_427 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_426 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_425 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_424 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_423 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_422 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_421 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_420 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_419 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_418 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_417 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_416 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_415 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_414 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_413 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_412 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_411 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_410 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_409 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_408 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_407 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_406 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_405 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_404 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_403 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_402 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_401 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_400 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_399 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_398 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_397 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_396 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_395 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_394 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_393 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_392 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_391 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_390 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_389 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_388 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_387 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_386 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_385 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_384 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_383 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_382 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_381 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_380 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_379 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_378 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_377 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_376 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_375 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_374 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_373 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_372 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_371 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_370 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_369 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_368 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_367 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_366 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_365 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_364 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_363 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_362 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_361 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_360 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_359 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_358 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_357 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_356 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_355 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_354 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_353 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_352 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_351 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_350 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_349 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_348 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_347 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_346 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_345 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_344 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_343 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_342 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_341 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_340 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_339 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_338 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_337 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_336 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_335 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_334 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_333 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_332 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_331 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_330 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_329 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_328 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_327 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_326 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_325 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_324 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_323 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_322 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_321 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_320 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_319 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_318 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_317 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_316 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_315 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_314 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_313 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_312 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_311 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_310 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_309 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_308 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_307 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_306 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_305 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_304 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_303 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_302 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_301 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_300 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_299 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_298 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_297 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_296 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_295 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_294 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_293 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_292 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_291 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_290 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_289 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_288 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_287 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_286 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_285 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_284 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_283 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_282 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_281 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_280 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_279 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_278 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_277 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_276 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_275 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_274 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_273 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_272 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_271 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_270 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_269 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_268 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_267 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_266 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_265 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_264 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_263 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_262 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_261 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_260 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_259 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_258 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_257 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_256 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_255 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_254 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_253 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_252 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_251 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_250 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_249 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_248 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_247 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_246 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_245 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_244 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_243 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_242 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_241 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_240 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_239 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_238 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_237 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_236 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_235 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_234 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_233 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_232 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_231 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_230 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_229 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_228 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_227 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_226 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_225 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_224 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_223 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_222 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_221 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_220 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_219 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_218 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_217 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_216 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_215 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_214 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_213 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_212 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_211 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_210 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_209 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_208 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_207 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_206 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_205 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_204 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_203 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_202 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_201 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_200 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_199 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_198 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_197 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_196 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_195 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_194 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_193 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_192 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_191 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_190 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_189 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_188 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_187 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_186 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_185 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_184 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_183 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_182 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_181 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_180 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_179 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_178 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_177 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_176 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_175 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_174 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_173 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_172 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_171 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_170 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_169 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_168 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_167 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_166 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_165 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_164 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_163 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_162 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_161 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_160 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_159 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_158 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_157 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_156 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_155 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_154 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_153 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_152 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_151 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_150 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_149 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_148 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_147 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_146 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_145 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_144 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_143 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_142 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_141 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_140 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_139 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_138 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_137 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_136 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_135 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_134 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_133 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_132 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_131 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_130 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_129 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_128 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_127 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_126 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_125 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_124 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_123 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_122 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_121 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_120 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_119 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_118 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_117 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_116 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_115 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_114 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_113 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_112 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_111 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_110 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_109 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_108 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_107 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_106 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_105 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_104 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_103 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_102 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_101 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_100 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_99 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_98 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_97 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_96 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_95 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_94 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_93 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_92 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_91 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_90 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_89 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_88 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_87 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_86 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_85 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_84 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_83 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_82 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_81 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_80 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_79 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_78 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_77 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_76 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_75 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_74 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_73 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_72 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_71 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_70 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_69 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_68 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_67 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_66 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_65 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_64 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_63 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_62 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_61 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_60 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_59 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_58 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_57 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_56 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_55 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_54 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_53 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_52 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_51 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_50 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_49 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_48 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_47 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_46 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_45 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_44 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_43 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_42 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_41 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_40 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_39 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_38 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_37 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_36 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_35 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_34 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_33 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_32 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_31 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_30 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_29 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_28 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_27 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_26 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_25 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_24 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_23 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_22 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_21 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_20 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_19 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_18 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_17 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_16 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_15 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_14 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_13 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_12 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_11 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_10 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_9 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_8 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_7 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_6 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_5 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_4 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_3 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_2 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X16_1 VDD VSS FILLCELL_X16 
Xxofiller_FILLCELL_X32_473 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_472 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_471 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_470 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_469 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_468 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_467 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_466 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_465 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_464 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_463 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_462 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_461 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_460 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_459 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_458 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_457 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_456 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_455 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_454 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_453 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_452 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_451 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_450 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_449 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_448 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_447 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_446 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_445 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_444 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_443 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_442 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_441 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_440 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_439 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_438 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_437 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_436 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_435 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_434 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_433 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_432 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_431 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_430 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_429 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_428 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_427 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_426 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_425 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_424 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_423 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_422 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_421 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_420 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_419 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_418 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_417 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_416 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_415 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_414 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_413 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_412 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_411 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_410 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_409 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_408 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_407 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_406 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_405 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_404 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_403 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_402 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_401 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_400 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_399 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_398 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_397 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_396 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_395 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_394 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_393 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_392 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_391 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_390 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_389 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_388 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_387 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_386 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_385 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_384 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_383 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_382 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_381 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_380 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_379 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_378 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_377 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_376 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_375 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_374 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_373 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_372 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_371 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_370 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_369 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_368 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_367 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_366 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_365 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_364 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_363 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_362 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_361 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_360 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_359 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_358 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_357 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_356 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_355 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_354 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_353 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_352 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_351 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_350 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_349 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_348 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_347 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_346 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_345 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_344 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_343 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_342 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_341 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_340 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_339 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_338 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_337 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_336 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_335 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_334 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_333 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_332 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_331 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_330 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_329 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_328 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_327 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_326 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_325 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_324 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_323 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_322 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_321 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_320 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_319 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_318 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_317 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_316 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_315 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_314 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_313 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_312 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_311 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_310 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_309 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_308 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_307 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_306 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_305 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_304 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_303 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_302 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_301 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_300 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_299 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_298 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_297 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_296 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_295 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_294 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_293 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_292 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_291 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_290 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_289 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_288 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_287 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_286 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_285 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_284 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_283 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_282 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_281 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_280 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_279 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_278 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_277 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_276 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_275 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_274 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_273 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_272 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_271 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_270 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_269 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_268 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_267 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_266 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_265 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_264 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_263 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_262 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_261 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_260 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_259 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_258 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_257 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_256 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_255 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_254 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_253 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_252 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_251 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_250 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_249 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_248 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_247 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_246 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_245 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_244 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_243 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_242 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_241 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_240 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_239 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_238 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_237 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_236 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_235 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_234 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_233 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_232 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_231 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_230 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_229 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_228 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_227 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_226 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_225 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_224 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_223 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_222 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_221 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_220 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_219 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_218 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_217 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_216 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_215 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_214 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_213 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_212 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_211 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_210 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_209 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_208 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_207 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_206 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_205 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_204 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_203 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_202 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_201 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_200 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_199 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_198 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_197 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_196 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_195 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_194 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_193 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_192 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_191 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_190 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_189 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_188 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_187 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_186 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_185 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_184 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_183 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_182 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_181 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_180 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_179 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_178 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_177 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_176 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_175 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_174 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_173 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_172 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_171 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_170 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_169 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_168 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_167 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_166 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_165 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_164 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_163 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_162 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_161 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_160 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_159 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_158 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_157 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_156 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_155 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_154 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_153 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_152 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_151 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_150 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_149 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_148 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_147 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_146 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_145 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_144 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_143 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_142 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_141 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_140 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_139 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_138 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_137 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_136 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_135 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_134 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_133 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_132 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_131 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_130 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_129 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_128 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_127 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_126 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_125 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_124 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_123 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_122 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_121 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_120 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_119 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_118 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_117 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_116 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_115 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_114 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_113 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_112 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_111 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_110 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_109 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_108 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_107 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_106 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_105 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_104 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_103 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_102 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_101 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_100 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_99 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_98 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_97 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_96 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_95 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_94 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_93 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_92 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_91 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_90 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_89 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_88 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_87 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_86 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_85 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_84 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_83 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_82 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_81 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_80 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_79 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_78 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_77 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_76 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_75 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_74 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_73 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_72 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_71 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_70 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_69 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_68 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_67 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_66 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_65 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_64 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_63 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_62 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_61 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_60 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_59 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_58 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_57 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_56 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_55 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_54 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_53 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_52 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_51 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_50 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_49 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_48 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_47 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_46 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_45 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_44 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_43 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_42 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_41 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_40 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_39 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_38 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_37 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_36 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_35 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_34 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_33 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_32 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_31 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_30 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_29 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_28 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_27 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_26 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_25 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_24 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_23 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_22 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_21 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_20 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_19 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_18 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_17 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_16 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_15 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_14 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_13 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_12 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_11 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_10 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_9 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_8 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_7 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_6 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_5 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_4 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_3 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_2 VDD VSS FILLCELL_X32 
Xxofiller_FILLCELL_X32_1 VDD VSS FILLCELL_X32 
XSPARE_PREFIX_NAME_0_19 VSS VSS SYNOPSYS_UNCONNECTED_683 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_18 VSS VSS SYNOPSYS_UNCONNECTED_682 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_17 VSS VSS SYNOPSYS_UNCONNECTED_681 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_16 VSS VSS SYNOPSYS_UNCONNECTED_680 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_15 VSS VSS SYNOPSYS_UNCONNECTED_679 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_14 VSS VSS SYNOPSYS_UNCONNECTED_678 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_13 VSS VSS SYNOPSYS_UNCONNECTED_677 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_12 VSS VSS SYNOPSYS_UNCONNECTED_676 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_11 VSS VSS SYNOPSYS_UNCONNECTED_675 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_10 VSS VSS SYNOPSYS_UNCONNECTED_674 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_9 VSS VSS SYNOPSYS_UNCONNECTED_673 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_8 VSS VSS SYNOPSYS_UNCONNECTED_672 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_7 VSS VSS SYNOPSYS_UNCONNECTED_671 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_6 VSS VSS SYNOPSYS_UNCONNECTED_670 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_5 VSS VSS SYNOPSYS_UNCONNECTED_669 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_4 VSS VSS SYNOPSYS_UNCONNECTED_668 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_3 VSS VSS SYNOPSYS_UNCONNECTED_667 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_2 VSS VSS SYNOPSYS_UNCONNECTED_666 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_1 VSS VSS SYNOPSYS_UNCONNECTED_665 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_0 VSS VSS SYNOPSYS_UNCONNECTED_664 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_19 VSS VSS SYNOPSYS_UNCONNECTED_663 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_18 VSS VSS SYNOPSYS_UNCONNECTED_662 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_17 VSS VSS SYNOPSYS_UNCONNECTED_661 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_16 VSS VSS SYNOPSYS_UNCONNECTED_660 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_15 VSS VSS SYNOPSYS_UNCONNECTED_659 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_14 VSS VSS SYNOPSYS_UNCONNECTED_658 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_13 VSS VSS SYNOPSYS_UNCONNECTED_657 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_12 VSS VSS SYNOPSYS_UNCONNECTED_656 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_11 VSS VSS SYNOPSYS_UNCONNECTED_655 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_10 VSS VSS SYNOPSYS_UNCONNECTED_654 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_9 VSS VSS SYNOPSYS_UNCONNECTED_653 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_8 VSS VSS SYNOPSYS_UNCONNECTED_652 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_7 VSS VSS SYNOPSYS_UNCONNECTED_651 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_6 VSS VSS SYNOPSYS_UNCONNECTED_650 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_5 VSS VSS SYNOPSYS_UNCONNECTED_649 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_4 VSS VSS SYNOPSYS_UNCONNECTED_648 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_3 VSS VSS SYNOPSYS_UNCONNECTED_647 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_2 VSS VSS SYNOPSYS_UNCONNECTED_646 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_1 VSS VSS SYNOPSYS_UNCONNECTED_645 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_0 VSS VSS SYNOPSYS_UNCONNECTED_644 VDD VSS NOR2_X4 
XU3 rstn n3 VDD VSS BUF_X2 
XU2 rstn n2 VDD VSS BUF_X1 
XU1 rstn n1 VDD VSS BUF_X2 
XCLKBUF_X3_G1B1I9 clk clk_G1B1I9 VDD VSS CLKBUF_X1 
Xu_gng_ctg clk n1 ce valid_out_ctg VDD VSS n3 n2 data_out_ctg[63] data_out_ctg[62] 
+ data_out_ctg[61] data_out_ctg[60] data_out_ctg[59] data_out_ctg[58] data_out_ctg[57] 
+ data_out_ctg[56] data_out_ctg[55] data_out_ctg[54] data_out_ctg[53] data_out_ctg[52] 
+ data_out_ctg[51] data_out_ctg[50] data_out_ctg[49] data_out_ctg[48] data_out_ctg[47] 
+ data_out_ctg[46] data_out_ctg[45] data_out_ctg[44] data_out_ctg[43] data_out_ctg[42] 
+ data_out_ctg[41] data_out_ctg[40] data_out_ctg[39] data_out_ctg[38] data_out_ctg[37] 
+ data_out_ctg[36] data_out_ctg[35] data_out_ctg[34] data_out_ctg[33] data_out_ctg[32] 
+ data_out_ctg[31] data_out_ctg[30] data_out_ctg[29] data_out_ctg[28] data_out_ctg[27] 
+ data_out_ctg[26] data_out_ctg[25] data_out_ctg[24] data_out_ctg[23] data_out_ctg[22] 
+ data_out_ctg[21] data_out_ctg[20] data_out_ctg[19] data_out_ctg[18] data_out_ctg[17] 
+ data_out_ctg[16] data_out_ctg[15] data_out_ctg[14] data_out_ctg[13] data_out_ctg[12] 
+ data_out_ctg[11] data_out_ctg[10] data_out_ctg[9] data_out_ctg[8] data_out_ctg[7] 
+ data_out_ctg[6] data_out_ctg[5] data_out_ctg[4] data_out_ctg[3] data_out_ctg[2] 
+ data_out_ctg[1] data_out_ctg[0] n1 rstn clk_G1B1I9 gng_ctg_45d000fffff005ff_fffcbfffd8000680_ffda350000fe95ff 
Xu_gng_interp clk n2 valid_out_ctg valid_out VDD VSS n3 n2 data_out[15] data_out[14] 
+ data_out[13] data_out[12] data_out[11] data_out[10] data_out[9] data_out[8] data_out[7] 
+ data_out[6] data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0] 
+ data_out_ctg[63] data_out_ctg[62] data_out_ctg[61] data_out_ctg[60] data_out_ctg[59] 
+ data_out_ctg[58] data_out_ctg[57] data_out_ctg[56] data_out_ctg[55] data_out_ctg[54] 
+ data_out_ctg[53] data_out_ctg[52] data_out_ctg[51] data_out_ctg[50] data_out_ctg[49] 
+ data_out_ctg[48] data_out_ctg[47] data_out_ctg[46] data_out_ctg[45] data_out_ctg[44] 
+ data_out_ctg[43] data_out_ctg[42] data_out_ctg[41] data_out_ctg[40] data_out_ctg[39] 
+ data_out_ctg[38] data_out_ctg[37] data_out_ctg[36] data_out_ctg[35] data_out_ctg[34] 
+ data_out_ctg[33] data_out_ctg[32] data_out_ctg[31] data_out_ctg[30] data_out_ctg[29] 
+ data_out_ctg[28] data_out_ctg[27] data_out_ctg[26] data_out_ctg[25] data_out_ctg[24] 
+ data_out_ctg[23] data_out_ctg[22] data_out_ctg[21] data_out_ctg[20] data_out_ctg[19] 
+ data_out_ctg[18] data_out_ctg[17] data_out_ctg[16] data_out_ctg[15] data_out_ctg[14] 
+ data_out_ctg[13] data_out_ctg[12] data_out_ctg[11] data_out_ctg[10] data_out_ctg[9] 
+ data_out_ctg[8] data_out_ctg[7] data_out_ctg[6] data_out_ctg[5] data_out_ctg[4] 
+ data_out_ctg[3] data_out_ctg[2] data_out_ctg[1] data_out_ctg[0] n1 clk_G1B1I9 gng_interp 
.ENDS

